`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
f8E1sXc0xBIeqHphsf3cJY5HaoqTo23wWTvYAfbq4PbGdbf3pqoeH8B1bRDMtDfh3GXrexdYE2Jc
EQxuqO6SCg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fRnF0s12nUC0Gu6ChqHa/q6b3kXe9Zy6M5DN1s53pMTcSkIHtk32R58ORE12IDaldqDbAdDvUwUV
PJnl+TlelcGuxtNawLmi+AcxA9xyAhXaym4nKcttp+iKxsxnA/7ruLlE5JQMdlvfUlJjL8J78Ltw
Dbkmmjg1UE1W0udDJf8=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mKxWBrU1YD5SxJA22o73EIfW8cmwKPdGdpNQt4NQClabAHu62zqZp0g+65Hy7wELci9s9oZCCrre
boHC3fwmxTgOtpvVfYyU9JNY5LfRdTp9TQdjV6TehSALBM6a5XCgF3diWI1k1Lk8NbI9up8iRRNr
+Rqs5xj4YOkGU0el+w75KHqwVDSm5g9S6ds9eMF7tc/R4UAzlgn552ZYsCIzUVnAGCHaDgm5K7be
3EkxIa4SPR45ZLF+pWAMfz5CLlx0FDdglZ3T91hPs9/qQnGh94TaTaHmXsD9dqSiVqxldt8Gtzrg
vDdIz0FRIoh+YtrFaX/AdIIBZ7md2/bMa8Bq4w==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oXy7169cPnrbCEF3oCShbXU4LCwsYzExef33f+pdex2KbYfq/4pckJ4ZeTLlag04HrvP3po8oOjW
plx+T05BG/wDyhKDM3j4a0nrizBlZf5D6mkZvNewx3zveTc3o0BQP/R+YJcBHyV/8R6CIqtwRhHJ
Q+22ne26AII78s5AW6BVF+u05ltLDvQXtCClhW4n1pzO6rgzL6JKraeDyHk5nkENVEgWphlaZKBL
EV5mhU1WphRC8oBaR9jXXUN25A8gPmebpJLzyGSTntDkThQa5JqcgRRLpHm75bfWZU2+ctT7Lh9D
3zYEyXKSA/B48KYxMyPa3Mtxsl7PGGxqJ+jpmA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
njXCaxI0ZrpeIsJHqmtppC+QoqLQTzoDBsaZJ1D90spl40rA2llUnGjjl1Tr0zYYMFK1f6TXs9q9
jNnMcWtkurdq+CZ7qRsXQ0yZWWV4SMqMyNoHCy2m21EIZxZRHnwHnm1cxBSDnUguhG7pjskygO/K
498ROj8T/Ke23+MxU3YFhNRQIfSWDDTwvu5+npW0Mhj6iz6wwh5ecCM5HS/95A9eAHG6m08r+/VH
ChLqbKbzzc3h1OVq1spLfmzhP5pqK+Pq699udky8u/zY7JV1Hdlkl/Gdy8N+Z7vDBreCXzp1mhhG
zhl3ioStjU2GilhQk7ZPB1qs/DFUrmMzwKtrvQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GJ5ELBTtiadRfLFYB1aBdbztJOGHP78n1I+Uj1MupFPJ0BSYP5JpWvJJu3pldWRvlrz8txpdJIQV
PNCrJmBDGQX+Jpg8FC9Fq9B5JqyfNSH1OTnLLuwO6eYgwexOT0UjcdwORX684j/i8FwskmXw18bq
4xDDPQwI3F3vyVOmV2E=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Sdms76Ale0JabjyT85uTFeFMThBxiSia9DPxOzJkQVFYDIxOn8H98YhyBy0+5NAWvuJgNUpwI9m4
G6vKW89pJgi1ULDyl+OZLHycgRlL05iKGZAOS/btTrNysliu3nbSmw8d15ZW6uJhOn59tYh11+Pc
/9vAQu+Xzux77/rjrOyCNWwEnTUaRR8HMztLSYaiPiU1aIbWyYyxTQvoYpnptlaz1umjCRc/rAsT
rurSnD9yhTNEfGxEc28HOpfRlQvrz3cu2Oqcmx19C5VomT6sD+Kbxrrl9everazsgimolYSLXM3C
hNCpDDPdDunhjCMlHMgIzwVQR84soZ41TkZZuQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 55424)
`protect data_block
Kg1cpuSdDOnL3knU5ux8pGUPAXMb7DJcfBmv8dwiR9CaP13cg+G9U6F5NwJBjOZPRxE1k7Kre+BI
HsKAzYNkOUG94By1wUlMUcvSPAPFy6EP3i4t12Q9O34g/2OBv4SD5lrl2kRLOBeG4XEKy45ELKMQ
bf01DnJEYDyJ8Oq1re1H6tJLZIaovRCHC2YDOW3EDlfxMnED/5XTe4Y8pvi1NRxGrCyttHsmSAWE
D/VZhAzeZCGXg1K7Suggt8Y94G9XuxdItjXw+hB+fSX/shsCxElXntxPT7qaPpqC+pCtM54DdY1N
uGby086b4bcUEuGE0FQL2xAKFJvP8ZTl/iclfSrnQnssLT5GkWx39B3Etc9Rvzq5KkngmWAUwhQG
ynbFdiBSqhhiI5q1tyUZ0l6CU/jEhdqmI1Q4IFeXl4Knl+Gj25p6DagPAeXfI/eZEB1T4F1MWRT6
xGzAt7APXCvAP91vTZ8ThxdEOnhYYpZ7DrsoGeJcBavi0IIA7tFGkIAtkg/1v8kVAxAN4j9Gi2n8
folxUH/tC9kAHvwJUD3td+ZudbDsHqT3PHbQEefuapIntHDkXxg1i7Uy/ls7qxxe2UasZ43bP139
/TQOpY6l70VR91H3kucBpdPnn0PP22mfBEaeEPflwaxw+WGDJXykNehSRkJvN5HHJxkAB2v7wrNo
Bc/yTVeo/Bzl+Ub1yYEsbJBr+NhcXZwoJl7jRORiul8uZdhsmi4/MHVsnqirBZvZcZ3w0bX+Pnbe
JNXIgnvRlL/9a0YXYaiMak9d/4IwMd/2cvHxclD1xYo2jmmU5qNXDn85ziK4MTh2wLKfo+khCNvA
q4FC0PyP+usAntBhowY/Rxk1uZVb3DKbT0B11KbQePsyf/EytYtZbXgUwalx4LENvJe5bcZKCFj7
W/hiKSwSg/AMEixccHKC4qLJNK1To1NV5ZgDe2T3WsPgvtjKq8QJy5+5XbmiVmqDWccSyMZopY2i
L4gXarZiYOaZ7fL0w/XwxagyNAN53Q4wJ/kI+abLC9kKLmqZr/+fTITQPa3LnrIoRSI3HQXdLyfU
kszXr4gHq9QTsbJDCV8NKjWnJEArz/lcMGwkgOwCLpQGmgGOA+rSO0T+yPk/JC7GQWH+wJOdG7Ux
Zx+998QnQQoX94LDPERxd4gKueIvlih2YkRjKoIowmZU0TBB9GBDu6z/KAb8IWE0ahfoD5s6vX/l
exp1XJB6YXXnXu9At9xpq98wr5xQNvmCagabnCjWMG9TlBiPaxHkW8ce12hiD+3z7FeP6Tss7ZEg
1A72HEePc/nCHeSOPKmfsqKi/Z87d18C4mRsLr5UMWAojiMjA4e2ssYhIbzjGH972jpMKqym1Tks
OVjEvIZM18Sh3JCXzbF10ZhEahOwbHF8Jre3DzCagSZy5ppvePVoEuqHHsogBKShMCgnyqIcoXaE
zrzSqMf5UOZePr5rhZmvVCSD3ncVUfTi/mxH1gjOZjzhvRH3rf6JKHky5jI+tQKzgvXPs87iOJ3U
74UD/KdYhNB1xu6S/QYYhOxqntMN9bErm5hD+XImVoXryloL1b07disTjqnCURb3lQFSXt9bavEc
sGlYJrub6WjlDAJBGNYjkOYeQb90KnIfIYAO2wiM+LIFpmV8OxA3g8VXbnte3vidDKb3QIr5EddZ
c0XOY1b6ujXMbItKvpn+X/IsNJYMU8H8U4vUVxhDjnfwx15z/nRbAjjbz/wAnxk6zPqy+S+Wff7E
3Rvfk3CisLFO3fT+Gq9xgE+zP7FN5f4pe6V0X7m18MTxA9VmXeVTg/Aq7J7PNgTVwQ4oS9P1ZYr0
c30yEisyjjINmY3Pf2SwPqzhGJLs7BcLqt2o190mPT2+qA14nCDR/6Ry7/CxuL6bF7AuCENAdZcB
JYC6Y2UFLc7TIsBMr0MVh41F3nDThLMAANsxo0XmY1I4gQwHOh7TSlT+8brNIScxL6yE9aLOWIhL
mnmF4RijH3T+GyrT6KrRuYWW3O/QIGvRlq5pKhB4aL/L18z5pFH+PeUB9g/Mze8M0/S0Mav5MyOS
mroog/+zKquXJGSUIoiIPumqxRLzWPKEGGLTglp9Gli8mPCdmU3moyLzRhpnAWZvpnmiKBrEM+bT
6ZX6NoHU4FiYii0YmJ2WxELIT3ufg+GhNihQaYviAUKgkNQ3JFsMDt2ZjmhCOCTnHOLCsHS7uBWY
NQ8C5EkE/VjR9cWYgtONB3eF5FrKXS7+5uO7uCPrDlZSV6E0bZN5ght1s6h/fLwwQBF7cRNVuL0x
VL2hdqJNwBL8RofgS/xUIGNxD0lXCxo7gUfYG3/sBxisFcGf6fuemTLIkTS/ZosYsLnuFsw4Je7Y
LlhbCy9HqeEapbwdJEJ92Mfl1dqIRKSPYnD0Y60XKnqrQL/sM5c/1uLxMxXz9woE64UQ7cD9ncMK
NFERwyOiwEbMPZvtr+VET01yVRA49GelaPA+rUhJg263ZOybRMotGJwYLiDI7KuUrdaMLx3et07L
7efA08Swm7blCO0wR9p5I0aG3cqF/vMUUnZeIiApielwoflIU+G93hgZUNs+KFHWpxPaKwWldgXm
MdTDkpc5Ic2/F+9I1yMPsd162qGaTsUwJUdbGS4+HGJmf1Pv3Abqn4W+HISHrSYULOHVE2SS9Lk5
xtimkNj6G+VbJe/qMMWpn/b8Ade7QO8y2jz2gF5SLR2fDd+9gdmIj7scsSDf+i3LaJH1i7Y/rZGb
WZ8K/2gqR8bCeNBNk/R/Vscck/98lZPJ1SGi8tNatziqqdwLoVhys2RX+at86RxEP7JmAEw3UFrE
+W7RNyD2rYdDweZ2TW3HqIO8+yDovyg5O9v3s8ExhPV2T59Uf7iv7lyI0oBA86s38S9v3TJzkyJV
LuoxMrrwmS+HzzcgZ8gv5cqcM0WKAML8/kcsWy8r7riPGSHZmnfEx1EtWTzvuoHUgRh14ykUg2DL
CWYvI5Tj/BrZTv+73qlyYaRCDpW5MDW5RxMtX59FqkXXmjKvH1MC2teOId5aBMEpNH4xHJAHrJe+
9DI/1xOKFbP1YesNVHFd5OOZ4ymxqhueX5sF2HYDyCRtAh2/KEx0npKs4qJz8tUnLv5etQKS9Al+
ygrnrOrj1KCPscojiHr1XHrm9cgZbW964qXCLIR+E/v4o7pl0OEmo6aM6kqt0a0gMP482C4Rape3
yCU/Xt4eOmz+y7n0Wr94S4dnlpUbicnmlpjFNLnN2r47/PvYQ9ypXW7YYz+7O6PFZFKft2wc9XPg
NJ8Kbr+QyOJLPBtgWbElBJm92DNL5UMSTzOFOw2kkitkKEPf4exKyVmSw4/mUIEl0zUAgPNnU/XG
Rev06mI1QIx00usHv5LjPOhiyZF5bYIbpiPHnMyJ/Yik3bg6vQoI5hFte6pX5VMYRi5KFoyJNQY4
OjumkMomPyGtJleRHGF3zU8v+35AwRgD/V361fcxZ0gwGDQ7mpaC8ay9yWe0CGU/59VomB471QEr
rX0hq/qRWUQQ8G1nB0rvpOobhP34rvEvN/0UgO+jfEJnNrlLYCLhjIdL0VeJdlW4E3fkHeX8Jt/A
pyNbseV+6JQMajV5MLhKW83wJqv7Dflmwmzn69GJTbzQFheCsnmgLmzeoW2/K8mxreiz0KLFSzlQ
S/aPUrgPCxLWfs+alACYo+gLSBCyHaYT4qZfcv5A3TornEANRSkWsFJTQ+hrmOjfx5g+LQEzM6g5
xFrFomiJ1zmfr2MRzGhZPE3PtsTNCbIfLBLOCknqsnJ/osKW4pkoIq9tK7lJvg+Acz/LrWY4bYcO
qeTde8b/O+f9yu8xdxxBiZSjRWhSTcyqOeJ5peOijaidvJ2odZYNxk8jOQwYMvt5NnAZjT3CC9g+
HCDNfoEt4YfQug5ZMFh0B0Q/x2SCbutnleRfTBWNSwCCGiX6wiNOoyJlNmU9g/llp0bk1TpZy8Bu
6k/B9aEug44CxfmST2teIz7iOCWKIp4zhfaQk3nRZD9Ty4X6WQsMfyDW6HeTC71JzBuT3xFFkbzq
+L/2ghc8Tw4B4Lr/eNzftCev7qAjRBVEZ83WRqE2JAeiX4Q7y80tHJ9ceESsOrMtO3DNVBbpCyqF
QTKSXv6Rc1uQiUgSWXbBAqsTcPhEKD5ng9+MxFTKrWNUODgBQzP0o69Mz0yuvZI7RrUncOalKEes
hfkWjwD0tRNNk4Lc3EeA6m8b7s6GlL/6bV82FGuGeHmUPR/dl4wvfzmi1NIofsJ4hKaXCD4giJ5R
2rMZnSM7IanDkK8l2llmnnG2hEr3MFDiK6JGwjizKytBVn62mzCIf99LI5MoP5sVbdmZl9SWd5Vv
nwnU5Yx6Xk9s14f1SFP2SrjBxlkvEUUWfvKdvSSFrtnCIUojTZBe3/7++IUo0AtdcwUxKs9ISusi
yKbsTQM4m1ZnRdLmvIKrN8Q2RJ/jnmpL7qZHAXJk9wcPTZa79oJ/WiYBb75sEOMIo8ZKcYdF7KBF
8GhDZ/xp30dxmFeGKie8IQcfXkr61TzI3ELIWkFDoskh3S4qj2GbQvY/gdV+4tJdKQDVggIRTfS+
hHwHxMRa5plZm3JjaOgWnPRa25B6y3XMsc3p7sYP/HVJrxiC9kfL9qTQPcYW0+4pqCC2TIVwAxF2
Id/ttpH7cN14BD9v+bTO5TVgPcaN2CDNJeGZ0zxdpTyEVtDDW+8Iny3KTJcTgMPc+bTosN3uKUNV
8zal5OxrnXAW8ANggQaxOZP7AkgkkQIRSF85Trttge6p3nQgrUY4CdQz+HCxojYEqYG64rkOhUaL
ikNr49zilo+Ivwx/GPmN0MXt5zWOPDtt3N1/tHQQHcP0Wp74VwiPvVh18ie+FlzK3+0QR/2b1i85
dP9tFo2uwpNmL6mXsN2pKGWwlb9X3m+sC8KcmM0+u0kcZi4R2etE4BCPqDB9GnODAJ/sW8Ph5Rxy
Ada5jt2bQb8t+XPjowu08T1EA6/okaR8evHRaZZoW4r2vSOCrGAm3XK7p2CRd91wFSmC17eWJ4pl
OmYEoqup1eI2DH8yiHQgap1f+v2SvR9oCEveXYxhyRK9/3ekr5+Fi13GV5DPpcrb2YURtJCeMdQA
T7s6WvC0i2aDu0y68/wR+LKJ2FOdlHgOMMeM1X7Sg7gwom4zt3bvHYF7a2geCG1bxILcakuzYmXe
qDZKbiUXKfevRrfctx4nQ786z/V85N2kkMfOAlJ0xd4+0FC3uUgxD+DqTEB2kOm2X7wJ1CFipwyc
7VqGOws1nepEuispyzGDnxwEkKi8EDES2wNxbMogdtyhxUv9KO/DcX48c9hQNtiSTCYkmZgHGGda
JaKcPvcW383sLQqBss3D8qLugTHRO1rgTVoK3o0f/pibRUsVbYxguCwN3fDJcZMLupxEIQyk2p7N
o9mM7TH47hj6xnNlh+rcPbLfNywQbgJ8mEAQGssGWt95ke5IdIralpaGP1F/PrQ+wDy2WfspzK04
/Frow0QVGTkt2Ip0B4YuC873sWalXD41j8H1WvXmIRUYXASKPQFJv/5y7Y7PzTrQ8L8fuivDLuYw
8F8MXaYZDFMPg1r5j7LcXatS4bf36bORuK7x/d3cP7E4+MMXMYfpU9DNIAWnR+ji1ANI231kmCLJ
EZBwNk4mNxALSQ1+VZXz8msw6RDk3riOdAMGYTerVuDqueiifmHZPs4aqMtRdquAeGf16InFrfav
e7KywbiyhaU/4e3s3bzUfZNhTbmHNdvZAwZ/aY4/WCenCVhD1xsEZPIuwh/5/o1wHIkw90Yro77N
clUxzbqTiGWQ6jFj4FQLFw1JlpeY1hh6cBPqK4CcUc3lMjWQZYYKtSSzm4SGOPwraRb5/Z/omDBA
l00DM8Dr+v1qxBB48WsvnfDve2wZfwe7WhA9AdnUSrhOdi4qr3AdwdS2aUb2w9bodW/cwx5214II
9dMIs8LO6VMKQF9GtJv3uf+8aqVWRdrx2yzauaMdgRO2X/AovALKLmq8FQN9V8DL9aWwY/FWtH82
RpjVN2eQ2N7UJ3oibbH4gScXEZN5VQ2jYuWK2Od9eMA+SHwbMrPafkzwJX6jS5I2iLY+CtKV9hSj
pzHc1iWUomcPyT8w929g2gFK9ZAHc/I9kyeg9k3eEeEtiozi13p5SF5kq+mJrantyrUxfqBxgJ8V
A5MzxGJmDdnKO7SzQLdgHYsMJeuCn24I01mQ87oBDdd2nCJhZrf6PHoC1CQfqhASbmzG8yFIQu9H
m0C7Aeu6qoTiIeXhapKCjzXz3J0rOiO5ITQH0+kEriMGr42E5GiMjZQnk5FPJwiMOD74UlPBJo00
W2mdECYaWFB0XSM1yunQgFyA4PaLtNNj0NJgq+WgZNYx9a5zxervqx41JkrBNSL4E8sE/gDH/cZ3
fFNnVm9TXgbFYTrC5UB1bmeUnGGFmLMdiKWMWnITlXXuBTsEn7soVDEQVzMYLgMSpA9S0dYGpFkF
DfSEvoiLZ/KwyuBY4PzGtLZL5SiPYd2mySo3Fkx7YH9mrq5Stp+xT/HWUfif9S2Q2oLgeAulFSWr
vyOqJgian+YurMnnLUJ8jW7yzFxssEuLanFTZDFJAatPnInhqh4txMJ1NqZF7g1HBKL5SAjB4RZz
Xfc6U1MOEkVVUDc9TBsXS3RUXV/djPrd3ieDIIABAiXD3QWu13VXAv4PqjqPyht+h5Js03lJETHH
ZnW2QPzNeQ4gZcjIVrYlWcA+P105XjMD0lnQZL8Yj1rhV6sgxn9bqQWmpXJ1ZI/2Mf7W18bgNUcw
Ln7MSqblMhzywnxqx+aFlXSpm8r58FmU3Uu6kJgNxpgPVsF9ZYlNORJhBL8pUJScK3jky1+hV1+W
nQF5NxX25BTYooodKoE5SwYVucicKJJo1VsdzO+oAMPGa4e2ZB18DqHzatTvNOBwqnLKpJKX6h6m
ksyxuPLX5Vbr1ozGusbcRv0s+4XyBHgl9yA+PdwWr+aUaVz45sLHWdBIBOLZ5Sj2ZTNI9e3dX492
rJwFNPGUn6bquJVlLr6XsMeNgxdIPYE3garw6xFszgqZStDBX+eYU3MhGpH0sHCRijSxs7HHiTSN
TH1bMSG34UjR0L+M+YdzRwbHZvlC+sHBqfhTlQszD2S8R/JsIBZvpAhNYQOM+xUDy/C6EHFSeNzc
IfYZFiTgzGj1vQL1bisB/ZMtWw+wyUnOMsYXcl1yHnVdJwQpUBkdZbpvvrG1wuTy6/MrSukWUYa5
za2CCpTU0zUhjedDV+DHVq2rFIvLEEnWK/Cd3JDqcCThin5iy2wjeIVabAC7+XasqPajFNlV7gNP
nAczOBhoMDDmxTjGEdrAnn3HhaKuCrm5yFvz0vIkuVyTOZjp9kq5T46CSNX44NFrCpyxnqKur25G
UtSzN7/Tt8LZ8ZNoBD6oEKmPHcVDRNbRkPfCarGbNoed/TrPNYNX0N3BCGcQr8aZLC8oqosKxxcX
pIah9KqCGN/JzzPq7fixTgQJvQWLjgveBmaTxgxrpL4NFnOx7GHlDoe4ZPEnkkaIHALUP2uq0VRW
L+D5CQ2tYFtwiQlUB9LYVul3ZQHmdy73oFHVmvD2DzCHho+ZO5+s0Q+pBFgTvgQPs8WRgQhDvnD0
mjMXOf3dDwLrjPE/U/uMgL5O992TwNf46M/1VIiaJb6yz2qpSkhjRyCTIpu3BhejE2+NLZTGNciS
df0FfJZ0GNbQpK6NHAeYD7KAtgwzbEDwT81SvGoAu+ya6pf8j2CUyoBEo+K4ecnEY0m004Xifocf
8RXBNdoBq0Dk7HBSM+QotV/q4SkQcaT2Qy5xuCyHwkg520nrOgqdAkyILrvFoSKxOfaiq/71sxst
YPx+KrbOYCE//tx4WDrYW3sF6/D2YIVS4tGwe7enlpJHcFHiHJrM5CycnQdJe7CkRe7Jv+7FCH2/
sQy9m8BzynNAA+7ipTE2xRfhiwWjjj4T+eYWucQZtvfh4utMmc+K3kkTDei+8TBCRSRfNRW+1+d4
TkY3dlYgYCRr7Kc5XKLyFw+P0eITQMBhrrI1L+31jQlU3uu4Wq25jOTKVtqMTDh1GXf6SuJjyptc
x6kkT4dr+FPolg05rQZDr+tEhiRiLp8RKD9LgkV3ggy0Q+DFf8m7Edf+IukwW/ulWgd/Seupl+Mf
WhPZcYWMlK2mUqsLj2bHSoDuMvDgA3x2wT5RFOqTVFhwbjgQlj9Q4TZ/sD2ga5Hzb5troT3J7oGj
ygkffLIk5Uv9epBecG+4q1DZkQZ8E99hi5clbrO9+KnIgKetvSdvwiIJWOa0nXDvR/FSdjIErdmO
klV/JIntvMrTkF2eCLZMQji1TauiaNfdfffK4TXbG5yorQCIVMourCeGfzCAYMwc2z9/D4rRegos
HRYY815dse0Fw0m/hRWUNvSw5macQCdbRlaTOJfLU9nvV615EGqYlg2xwhTrbx2AtMhcjVdecXa3
d6J+elUfF9wDLnaxPRllxpTPBAz2sQEvc8PxixLIdsMdJtG3+APWIShfK1NJ6fO1hSoQkw3qWL5W
7PDq+6EOvpot/QPAxlhLPL4Aj4/YvKS/3i1415GeQGOiWobL0LRJMQu2qTMZgfRGucFzdfgpljHV
6quf6qxrEvfv06jnUqrZhyQwT4YNP+zSSGa/cGy48/BTJM9x2qVhQw31DRI7DwWrbV6I5y9avyrc
WGyjK8XtILhAspneSIf/xsK8iKqdpD8Oq5niZo+fZtOTbfrg6TJ8b2ZCXxfhmBcHtD1coqsjhH0K
PTlajGCFFGNVx87Dudg4z0/Q/FnVV8S8fTvKiYwggkCHnylI+91052FKebLe0NFE0PWUPuhIhaGx
V5crNX/E8XUZNaLQUpN3nq3cxqX2wIwRrA9T6ps8tgmcUT2Jn9mTddGcxXFhZCyHAPDh0Ks4laJh
QPdTp2QRXoy56DljKlXxfinfnbngLt0V7n5JnNwIutqu5HuYpbpZGeElnUUBAClRUbzWqyj9cCm2
z92qC/ajAUqheqR2Q1dmhY9IyJO9r/O0vo2m1n5MdU3rAL1PjhimCbdSIdxRSIb5aldnUp3bQfB9
YhgAh403d1uEnwAWzlcTOLTFrZJOeWt1klnKRrGYHW4e8j59Ig2xYjxcTSlJBu3PaMp8dJ7U3RBu
LGgfwJCN7oPqxEZSTHvWKBpku69lLO3/gkqEeSD5+EIj4vtP+QJmwEgWLe04IZE1w0D+meQz7TzJ
oCkXifsPMw9FCqyD4ZiMAF3AvuS+AfitgCP4q0Gj+YGe/ITm/wod7/0RZyps2Nqv9Jv8hTp+3UsS
dBoxxyx69hNqzNNlObgWwCZPURdavcrf53w/AlUI30/T9lETbCWULMsjZ9veQmxxGcFgELZeQrlp
qkXxsXajxHBjV3830MmHnqItP/5uv4bELHfWYtVhlc/0j7SgrigvBhPkCfdeOzldhOvbEouGsDwF
O0ZDW/XVWGW+rhAPkY9M3KPbdWAfTJGAhBvWb1je3yYG9qTqhGkW5/F1irSaTTDk6tL3tamxnNCb
My9rvMRsnkNCXMdgHo89D/HZQdSkSlm6Aqpx8bWTxd6u7l7PkrrgiXH9ahKzfRKyki7nlcPZUzq4
CbemIqMsE6fI43whpWJyLS6hk1SvJ+pHjxbtVm7ayOGCNux5MaNv46tdFkURam2whQWiDTmXhS4r
MXifwLaFzMEYwo02eQax5jroWlNqwRJyZ1X+LGqZryih+1NQH1DxAr3pbSFmuXQDyIph1UoRJFaN
l/3sWgH8/q/PoOLYgLt6hgCGLEokuyUNuK3z2uPXHI+xaDjuhcRFAGNp4+V1K/uf8C3aYbko/pOD
dvFM0TXfnMpiggsPW+1RM7XGy8ss3WvaX78Dwfo20HprhVcyV9zMGkM3XiqAdSH5cLX9rfdJTY1t
MlyjYU7wNzB6xFXZN66kHAHkRbx1+q/La5B0xqd+7q4P6haZlyUn6GdMzJ9/4tCUBpcg/AtJzQeL
NwqXspmqFRPgZnc+HmNPtMBs3PlQjVre5uh36o9ZxakAxn05wrCcGxDUhmrsXs/uDZ9OV8EBBxY4
QjnsOLprUn6S4GxyqH9zr9Cp1iUFkeTtFUp46RVkQz5lyPYuOrTjSCtSjy6FoYU1RfY0MXJVNDIt
YBwDp6dQOJ/G+k30K+5K0Rb9vO1JpesP81H2oZyUJzWptSV84DC/XUoLJAA3bXxQRSF9mxh/X6SP
2RhiWdaQgW7o2qiyzCFpCZ8r2oiffk6xKb0IQcYnstwV8NXUPM/G9i5kVIoqdXUt+2/pDJD9LlBN
tyXd2EMl6sdHpWUvp/nTARlVLDO3azT+smTC/or9WGomGkUtyCKDJ1Yz4WhaSmhn6egg/c6AJTQp
5wnq2i0L67gAhU/O3hzDkdgCZbSDb8+kyC7QhrsNgxHc9Toao2QOby9QLF2qCZdstZfA9mXDj/Eo
qk1o3MdnXzSAz0y5HyNLKt1YOMzvmQnWFcHfPnFFx/feV9hLXlRHy4AzXaRaK5WbH2rnslsR451E
wHdbhKC3NRqFtH44U6bHpII+7vLeoze7r2t7f1FJT76NxZMDvP7WOG/0shupDc56Qs1AqJee9TDq
IraK4+OwJWQpvIhaWQ/3FQEAoQ32YFsn0rtwfMAmLKqzxS/6gIqORyZy8kjQOUy4PCcZoLeEZpvd
XfnWbYcMlZv4U7DpiM1aBuG9HZl/nSR3aYWvaC1n9NB4EDB38PAiyKqzgfj5E3Nc1on3lgrNF9Zl
up+jb9/sC7JQMKBXK3YZu744u4NiNwEhAkDRjidK9Ojh7KDbzfqnSFAWhi8Op16lCGhyW31fejoV
3ki52zBKIyq7YfytI394VshqkfrvzCJZLTTkzeY4ztWAkj7LXqq2Em7PGU3bH3xT2fRmnXKREbAk
lLMGtKT620GeM/hvE/7MtwOQXg4ggfo5vh2uoDUoaUsyDe3bfs8thxSzYDgAJMVURWd7DXDWGWt/
JsfY3xlpq526EimUlOdIIlknQstjFk9zjKlkwTx/4tWnmPxDEb9SmoQ03x1+j84+2Y7tcTtBVF3A
XQB6WSV9q1OBN71x2F0ZWMPDayGsxC1ADcCDs/phb8tmMJq7nYUqC8KjE7H3T2oSIBq4ivjIlnv/
2lEyKOQozqtGFFvdWAdief1O3q+jVRi6VVe9Ge1DU8fR54lYvFWHN/GoG1JjRuJyLoWPWN8oFfnX
OIhToyGZsSaEzT+q8wfdOiLWm+/Z08MJmEX0qqLdCsP3gPZHAJqJpibQZkEVanD3HjVgvbTp1+oM
lla+k2n04HbGO73sDTbBOOV/W/sLGLCplmxTsfV+u+ElWNwLZ8SdaSKt8R3xbLJ0XIM2yMZK796u
WSivx4ytPR/mea/byvlIgtgZuab+7N4Zk+OS7i8l2xu+oM7W6XkO0JTN4aEkUDMPLGLs4zYNT5a0
J2aOTXFSKlv6YZty3+r8tkKP+77F9W288oLQunhLE6zDNwq02ZjLUYOYxkjwPyEKHSqt9QTQqqI7
vRD8pr7kXo0JRJEttevyJH9eJ/Y5AktVF0k8pTPx5DRluAl7heU9xtRjn5EqlA4MgRodUrDtHfXf
k/3NY+NeiCxT8nbz3krfvx//N6PG6W81k12gZIIobDS79NQ/ekT7pe2gXSzkdbLWP16mtcbAdW9G
NiHXtKPw+5lQq5qbqEWqlhugmRyLjK9cct3iAu4iDrzFC/+14Pes+kidmbpuS1wyMCkpEuCpHVWR
ETwKUYblxyJAQDfn91xyJsKYo70TSgaTq10ijy3nF+L/v8QIzhV5ZIe+CWCrv1dMEfnEAgPAmm9P
JgdVYDIlZMOzXVifKziYuWpzZKl7n4MkHlqE43PvxPTMwv67gMqZ41KdgeKpFdo6tmqj99fEE9J6
E5GZ4GPc+ZGtr03BZ85thvq5ocSF8H7FFEQW76WeAyxjEGGQFIMW5ITSOWS/NvsK35waH2je1nvn
tY4JS5KhPLG9GcKuSSXJ9CQwr8ZKIuYbqpU7yj//QoREDFzPUOTZry4zRVmyT1xFpjIygt5Kc7IH
5L8yKCqKXFffxF6HvI0fLvqbSnUHO3gmlewqGFCDrBch+IDlNOXFnBvboulSLv/t+6euEHV7cXEu
KOMqNX9QeShfyrj6L/y+wA4EDJsOulsxk6ZZdISbuCFkb4YepDSzXNsbsHZ0uKC0iFk9DvD6MCff
+Cccc10fSHX3DzVn7TfLq0h0F/1ElRSpoL2HrcYi7+xxYFXmY6UQh/73iih13Ed0X9RHZgzNKBk7
kyVSA+w3AQga2mqVaQ3HLdF5w4yG1jsJ7P2KpKGqW+K9DcSHYHhZMHA9PA/smIe/KnF+s1XZdJiW
JQ9DahXa/kz3SreVVyFUOUxi602p4DKqCURcI7HbDP/snnwy1xeNqIJD4q3rmUayyu4ns3GU4d+j
9j0CnKpgeosNQ37he4W2rADWQ0eHaV7rGgcZwIFexWS+/GE851lwGRBSZBTCyDLv3OM/kg5+aIW1
Yk2egCzuxXgFVzaa9sLWvgZN7CFVrLqURDqepuwGRvKKtlrivGfbCpijx1oMmXn/i3HcEgxwLbw0
FHIOKm/pbQ9IRmRiURttvPWpy7beDeLXZtP1GsJxcPQ9UmcjD1F37ERSusMYyDW0YGeZlyf3Fkjj
rSwZq3bSkUBRFSoCDNQCu3ADDljD1fKnTrIMyvq7K9XiUjtqRR/EAwrtM4Ika6CRlnYj0jwMD+iA
eLXsFvl/rz5/q9xDX61yPx/cWrzH4EWw+WSXThB2fDlP7cn58tgL2giqS16vAUAtkl9z//5b69Sf
Nk1pydU/cOrJI0ODsXrm69aHwyQ2WQrq7nyQOGlZ35hmfOEEu+nsJ+ELf5zOuT6UVJQvNG/A1mRp
L0SqBOu2XskX8WVLu5BQWbJrHAeFG6qplISzoh3XR0ckUc54mGjkFceSZxOVydWAGH6Y28lkZtEA
hO17oEZv086LsYAhBJB/4e3l2/q7W81CSMtXYIxdy/J6qIrXHwq5mI8guTVGU5s6Hlfx+TW8pLp1
e/wV7PfGF6kDH1dVUHmYo7zq6Y7v/bohTtr5R7tsfG+/5PjCqRdXChXoRqG0fPx2r/zRe08BGrLZ
iXbilkESTySHhCJ/Hgp65SNKSuczqJDNOrB02iHATTDWKn5AUcZ6ZmzyXEXUH+2O4qbE1Yz5pOWF
8oPsvtSEi6RmCnSOcp1cUiwndxvt1FWYtRxbXl0vmagbH1fEHkUK/S8YXoOcurzdwM+alRQYfXHt
c72h+EkasoKlO9tcs1c5jUTrvxlqU0XgkC7Qk+fhCx5jU5UOtaGzoDcKLBxmOI4aF12nGc8bwAsD
IwAHzVH98Jx7kxj7Fy6PfgJ8ffjj3XjC3RyFr8Pnu2omHBEPEDiyk/IQkYvOwkfkSeFZy29RlZMu
43Kw0PvU9yjiCG9Wu90kHfjSO0SzC+WxD1WpLOgr9PZ0i7B+Z8UCLFxSB8oH2XzoEG+8u8pQEhOv
2riZr3XW/bLgoG3zxZ+d3zYkUE173KjdKnjqwtJsidRHc125hWL4YVHSCpQW0a99nFb4rdB3X5JT
5xcqoy3CP3luSxT6pCSRnToMArx1WIZjthemZhxJBsX0NUmXZpOkOuY8e9uc2ZRnjOGmI68mYM+s
OkXgCc44EIqGsGVgqT7lCohrMKaXFxZTtTj6mHqaqd1kMSzH3keUt7XUFOHrIbmqi2RGxGXTvVbX
xW5qCARnQF+/VllcSnzZm6U8lrtBD3Esi1T5swt6hRMxLOsN+qYKjjGIYpair+UFeJiLMDZZN+lr
jpTxc4lNsdWr619+7n4YYOGq9qRbzEDWizbbLwiaGYuU0i+9bTjocdGK0UXEuFNLBT7DY6H4cFyC
n+0PDuLBL76rz6UaXzC5QBfIuM8RjGa8nCmkKXECDVBSIftr00R0IG9qTqfmJ+AKQZktcZURYDLM
CJPBGsrZWJ+PTvjYWrGUp8EXP4EqsQEG/Qq0K7fBUbks0s1dww5YVjLdi8nHrFkuxZbfC8IhB+cO
Zb53AdPA+gN6awHG8VV21W+vAB96wpYHXo1dTgL9SGZyaG/j+fdrx9LKQ7XrfqILRZASAS6Mngyc
LvXbjdtFFB5bxozSmHkdF0/BhMRnpUGDr8H4tHX/VGsIZ2K6LLWapnz9kMR6B2Gb603Zb8RhsOcX
AglWSdd3bCu5j6qv/GNtr2cff0auwI0T5t/1DXZaDuXG2j+8QKZDfh3mh3xXj+y0pYgx8Xkbb7X/
feG/vhLF8FrQaufpzmPPapm/evwXDHgeh9gi85ytxRTYaaZw572YwOz7pKn887Hb9jxjVl3K2g06
O2eAs9/Esa7jBkFA5XnezGHFSJ3lYnsjiXxgkbhfVywhCEIRRmnTf6V9lg/jNdryOtsLHR7aJ/y/
IbRrozFV9mRG7dVFaZBQ9VrKfpGfbqef5iXL8PCi/fsCp7t5M5OwJazJ1J6ccyBLLw+JmIpjmWHz
PzUAyu+SfACZgBKf6QkAAo8/PatXSjSYr24tlIm1fChsfUfrV2Ylh1IzCtI1QTB1j6xqSk9VVL9U
LL6cdyR7PSWxBrOUSKpflXAJzheS6GCAXtmKTfmJW/fo8NMr3FcCBjWUyPSYcoYSRsGaAFJ3eZSc
0CQe35GdlnvltfXc6wBQ/1+/X/05WSuvfB/LAgDOWxOt5dxswFiJim2EpkDygL58oyaq1uowLlE4
F+pohzFrpFMg0SNUCksL49ytchuGpLBNmvNZLNtTjvEzUbbAb/wji9yoXYVXeHJrNhvGivtUdAOL
t3a+OvcXfh5vNxm8CHVY0tLhezQ/AshaOJKGipHl2L/wXAF/AMxf590uyKJ8P6neWvEGXh4E2YYH
PLa1+J22pcmZZ17Pp6ahDND4MWxjWOT4aL6fmoesnzFf602ghSd8Wif2WyYvkXOyt2THjtRXbnwC
Ft2oBu8pKByNGNAYdhywKJU+0TwcPph069UftA/9UCRYp18rG0ZmsMWsrBsLKkXF5Er5ooM1k2zs
ajAqu57ZBhzrr3xI3fGmU+QNUIUGd2f+4eWiiFh3VHKssS1wnNDqM9XyTZEk/92wbe5OMcS/ys7b
DOco9bMV+CpgUEZrDk7pAHuegdjCu/bmTEfiAF4EW03owi5ny2aVcPTdGJLZ1yifmsY3nBgiTd1K
/ZxamtypVj0YMryem6c84APVvWFgEAA24SvufDmunmMDLI3UTuBnBs+36aJUl0dp4NHZSJEal2hC
IGOX1a6nNEJttjaWFzujkYkOiTeSZ9F1b7p3dJBfWu94Qca/UrwJlqDNC8Ce8ndC7fDZkHoXKc4a
LtI0Ge/7WouueE/kAd2XpqnxDVjSCMnslkdXLDko+AVEDsEzkgzzg2yJFoN6hEdiW6D5AA4pBjN0
RuATYTFFgMaIUPLbY65xkPtG6Hyha3znoNowY0DYHQm31FlQaS0OAM/eQiBVnNpzBt0x+DVduH2i
7MY3rD3KPQ2TADY/EFyaMD17OxtgM9BvaG/6icdwSrDwC2/b7r2VWhRTKV45v912XqLhGhEYyeYt
/HPT9GPq7scPp5qpS/dk5+8j7cCMeofvO39e8EQF72vEAwKEFc4X5FqGblAW4U4GdvvVpSHRHrEX
AYDmtJkrmbigxwK0hDnyvW2Bfni08fJor4dXVImqg65iOq+rwCftqvS9g7SqGafGnJEmCzsW/O94
y4JFgRQsW7FTFpmxkjv5A76Jzia3mLuosvKGHjhWPgHooWWLQnCUXP/hCiV5bknt8+yQbNifmMij
oKyTt149I/HRIKB0qHq+t+mnY3d39oYnEidCKVyxkGxsQqNnCjxrsfKpUrskrwAZkppMOLbikkbi
eVcKrV1tq2cFsgyF0qOa84A3Um5BKLA+bVIN/45Osm2BhrROVkSVMktygmbCy+/5ca3H/0IYcCuN
b76ju9GnNdQbuKZg1uiVaqVxt6dlbHDV9/Li/eHIS7cgHGugcw5/749wH7V2d3oCAnqw/6z2z1Wc
ASmOkhkOru5jKuaraR9SEqNcR45/Xw0ITPP4HDAMssDVEbXgIXi/OcTRtA7ZgWG5Diu5uc3pC4mr
xRVeS0Ua1OMlXQJK0G55IF1YAOEzQRXNTF8C8IFhQwR6eta6YwIaYL3Lw3+rqmS3qXCXyzUkHM5P
G6zFmjx7oDgwYzKC+LG61WphYCJhJ9uATm80AjhMgKqYLy+CvxMG5ipeBOBeCelCvBv9Q4B6ht7S
H8H8rbFXIMTSrk5qt6HT9jv5grza8IZ2N6kHNSqKwiN9imbRbQwMpEtoqR+rAVAqEXwaWLHEcox2
QySG7M3c+z7+qGy4v5LCw8tY+1brvHR+jiV6lUssuEw0Q873k/JVJpTd5NTQZ2X8TQiZYTrFSs/o
EpIiI3KbJgq7IXBVd7DwSoLgs4qYGZCX0XhCajKvgEDFh8erZRXjekd1hiVfl3w9xbXj//AN3HiR
tuuj7nZ5vinesXAEn9m0aCo14KROAylKi83SjBeC+ueHCnHBqyikWy/IJc6gBnlZ7O/Leobef+x/
kMVH/eff5HY/MXfa//QzlWnS88f2w93qIm0W0CDO0grDZ9Ui43VDbB6kIEhfZ40E5yr5126NzIKz
C1ChSCdaYYOnFbR9SjpUOXb5AOvoqavpJIeq/4EmYvi3aLyjDaC6GYMG1IzyPCKxlpvzmcDq/ohi
yxZ4q3Vw52v8loM7SJfYUFz7ENe2/rpaBjO5/WfPwKy+RITyan5TMGFZiduWkVssDtBpigOn2sHh
aCtVdWA8en+7seqtlCJszS34Kmzw30SG5k+vU2hC0hJrzDrnFaGK2yLYJO6RHavlU2KwkRPF91+7
WtBkm9Ak+TgJ7At1L7A2FUVpZ7Yh9Boj2UR3CgcyJDYPC8+S2euvEBxiPH3GGSSxBWcPXHgFa4Ns
HmC+WbEu+omXdhiJDigJc2b7wBbPKglLgkprC67tKoPybG/zY669C2ZmKDR8Q7Dpwa9T93CS/rln
OEvEAbsjjfypT7/U7eMmwQgtcZD5EQC83AeuixboFDh37c1kVeTGIsDVjvw77Vg7yGaIui3GZLTv
AcosKWdpayNhQMHV+KvBBl1wOB8ioKP0aGn9WDpqbZcAS4dtzBIABZ1mneipbOvgOLrDtzxFRGUK
hPWss4Qi3IoDZ+TJzcsC7sDQyjqUo0QJdP6hJDM8jZ0t7XNzxERNGvvJdVVQ24qi2CfAgmwxv5yO
p/jWAJuieffhj6z0DC8v2sYBzlDsYKuU1oobCLa/3gO2Cfhw6MlWGijpedrRlVe6r67HR9pYznMe
K15SS0a7OmDwqmpbn6rr4dEG43niYLl0USaTp+Vx481a5sQ+mLHLkY0u/UV53RK3fuUP7K4cgfG2
6lCbOEymcLm20zvaqdKIaUOePAESJYRqgRxwjb68t29bOhYUeSBGAMGo+QUyI4kZD6KsynhxWjSh
5U5Da50oHBXApT75tTE10fiVC1Nv11VFwpz+A+b/Q7lK/2S615esRFWWOaBM3jZjaE7yFZMIQVCF
oUfa2iQaznqh3Zy04WVutMa3rDCvLPN2R0KDtNPhOJcWvv0AcE5v8Xne3IZYkHPTXB2idyNAiTm3
EYFLCnvkol/Fg0QKNSnipQu5kT85jINWeZKKAX2ZO/aIQpKz9DiSXQE7aA5i0wt7Ko5EZpqKJ/1k
uXhjy9JXS3XpdqJlGDT49/6sDZMoRxUvJuCEQ+Fe2IC5X9k1s0hLAcqcmcT+KgC60gmocAV+vFqI
j2lrK97gIckiUNq4Q82oXlSQI/ZSOgLg6Ie74Ks5AeSEUCDEQ9WkIUiqjiF4mMXc6uIa6hKAOHEB
TAzUf2YA1uz5tN3M7ow+f9JntN2CydIFU/KQ+FYJRGQeZ2V/HMvDOiQzAxYSGi9Qs8hticNAKyov
sOTK+3tVxayLLWcofA7G/5BiHim8vc0xlEf8qjZ9DVe6q5GJqkHZeLMhMFf6yKZSSVSThJrVv6+V
/Dy7WpCPxNQlUZrMpw+C8mfTPqgj4qAXr5fY3sM3M4/enbad6Fqfqb1uVUPKfdW7AOQlNvT9eH5d
k2tgaioYYhpA38fo9mUOM0xWcAdvP5JX6/3ZdUkHkaCncaA7G6EuTQ7aEmYiPYRlM8JQFhxkAJBg
EVuYXx0Sf+U9rtJft/aUQnjKz2RYRp06qr9SzFudikETTrl5LRZfM+xk6npcwr1KriR8a6Rwv/PH
12HtRCK7F4Yg7d8ajyVo50mhft0R5F8nu0SIAuQ+Q68iaQz32znwX7NsuyjltsBBQMvIt2MhumIF
00Gi5ufuHd/nkCn/MAyA8vXC4dP1uxX//bwKxGyWnR8dCf4pcPPRR1gZ/a0OZgeeqqMEGc2p+onz
0C+93IaO2iR1hMXplvprddndESjy4lnd6DJHiqDNW00phLD9nkjhfQRMnhLrkThrciCMkyoTFf8c
qjaWC9cpHQC5oQgPAXYiWKnhVOFIvBC4KyOTQogWyO4vFIkBephigr2vI3pB+6s8lJtKpJG/fgFp
DC8n856I7KI0tWSmlXNMUdjVVPMzuZFSEf89pDF+icLy/htPd3CV10EBoAyy+jdWC07m9la7AWrx
P6vE1JgRxx8T9CTsg9MOdVgHE6oqLN9BciGvdbXSgXfhOCdJAmS4DdabcNDibzwADkjVHfn182ZU
3Byu/EmPhzVFqwS2XaiuptwhcFiYep9A8idyBpCGBq9jmaaNNp8C5/LU3BBYTsRz6XG6u8ddnJza
YKGCIjuw2Jwo8EsQWi95Mj5z+YWLS5XIMG40oGOjeZGRq1U8iBNytU4hePz7DfxrdWWN3Jfk8z6N
+ORqhJXdFi4FZq4wmAntbTxs/HYO0Huj4uzIwhT+2N2PtyRjWOMb5paQm84B4rDmijuXXF7JHx7l
ZtAkuR+tbwCcZLwcfACny/PN+RiYc2WzEqjKrdkBzr8zFOvUnx5n9Zc8DhMhY/JgZqXlVdGQ2R0z
aE/TsoLbIeE2Scb9aVkvQFfGitQy1qHYNfVCvDcbJ0K/X9W1ncNqgdrjQI3T/NGxh39EuQEKakXH
B8pt8prz3HS9XeTpveyhA7N/emQX13tODIeu5v26UC2SRMbTqpkhQO8ntoauHNzFYryAlobKoMOJ
aRBdhdh0X+adjxsF5DSInubv8gWoIejPD7gWbVQ0qgKYaynClNluciqwIP7E06c2oZ0mx5Mmr3iS
mA/LpAT+zKy5yiCP+ABTCTOT7rru+repvAB0x+BFKVgdAQB0KQ5FinKMEbtzKH2HysEgbhDT7mzV
pdRbRYEe9shtiTpTJSrgliIlau9Psa+vq3SGHD0TNLVa+tM9D1Iy8b+xU4qobjbCqE5IsPu4uIMl
W1t38OHZvxwfTm6OJT25ptwLGxteT9Og5jFS+w5vNz+S3H0xKf3wV2/mw/jn2ui0/qj9FdElwz1E
v0zn40jgWX3KvTNPrLXH1oMSDfY87UaUSOeS5Z3RBc+OKPfgv2/NIlC2aB0UyhiPRghXfeIvCxTv
mzHcJpxAvy4wMpdXCaI7Xxf83cjJK6sSkIXDI5Os9oxyxtMpjNI+m2ju5q8zQ05yn9w0MghU4GNL
Ry18P+3qAuQ1O+WYJLSQvPG6sBkoGUcdXBjkK5i5wE5w83P4CyQ/w49kyIAAVCREZ9G/rdVNQIjW
50uhSq+rUyKrQo57QPHmaIQpJzt8II1uKMl3aIkJnNkwgduLSUiKBicPk6XOs9b4kW9PaBEgrTxJ
6sf8EKwHIgSDT/LJ7JKzW6d6t7PEe+x7RVak38RIIyu+LcvSdRQPEkGCP5CnRjP/w6u8RGIwjnz5
+UPWI0yxx27krtqf2n1+f/ge3b1ZZJlPJ90awIOV8RFfi9SaTeJ/+ifiq6STnDOBGGsTqDWgfOsy
WCRVHmY7iORBF9nrpFmE/UgTbhY3f2V5mvayzWjQDA4vGKEcxw/Mk7qIppfR0MhkmW/CBUL/Y471
HvNXZNcLGDk1SOsUDbxaFa8EB+aflPh700QLq+Q8xi8LbFWJQpG8V0rTRis+oPQxZ6nnLFO4dEvH
FYAhFhydk1fuaX4RBnpYYd1Np6IrDTUA4pt3uLQkklUj7KtNGjCqhF52PdgyKg2hqiXSMoatPr4r
qphJug8QROhKOuMy2UWiouLBw/k9F8gvtHx6tvBcVnM2/qIRIBg3L/P/V6DStvMG+NG/sBazBI6w
+rk3aHDAFlsAHjSZ6J5PbNf0crMZsM24A8+tutThfJMAt5flktjtjkY9A5FOsQGoIy6nates/H64
RQ0r9Nagqgc2ypIytd3Szsk4e2wcCSJi0cXC5x4ub+yvHSA3QHO1o2E3N5BA7fJQ3FD2nVwtNFRt
bf42KbEW+Dgf5gMw/JWEGXAY5ZuArfviiF2R8Ek1vleEfq5tS4VXEzqHAuYmRAKzLDLpHwWBOp2S
Rck8kYpxl+muR7XX3Ad0+8KlWMK1iIua+YHUebCvbXzpcW9GF2ZAJwuAtbOynhfwxA2C/+MkUUDl
8RY8nBxCA+T7ujVIHChCzdohA1/WwFSjlL5Dg/e7fDSZBuv2vOuOSaVxkvbjC89TQSsSO3CnVmSK
t7GraVP+sOHBXCrPVi7VeLJ7sJb24YE9vNPHf848BPQefNv4of6zVpmxg9YfAqXkVHcODppPCRtC
7mUhn0utR+Cuorlq3ZkiAzZyIVLgDZTYLxB7b7S6LEwtBhrBAyw+3/PLzVRdnhI+SDXjfZx1zi2i
p4WUxYFyhtiGto272cvTbxkJ/qpYrJ46KxDvagL0DZJlfsfJugRjOxG8JYmqVNiqgooyLSd/LZoM
tEmY7XXE7Vk1h5NIY69Wf8Za7u8HsA6eK5wlukpDWXZvC5ZHKrHuchfLc81fzCNtg0x1pF8pNBpk
17zy1lhbX/XaDzHTkDxZ2MPLaz52A2Ukf2vc+c38PDMa5Y0hFg8Q2G4KK8MoC5R4HLsjqr9kGFLT
GpZc6OD52AQLdzlsUoNKWlCd9o4sFOHdMpGKNOM78VijrCk3+Kgmq/2Ew3o74WW+bOiMWSW6MU93
BC5SBstKLleRdZ4W8phutkyI/QC7+qhRCAdEqX62ZoRQlYwVS6pnVJPfzPYvOWjA/S8KA+OA0a8D
NyklwFyGdOGCJFExnMqMpOID6oYWGL+WIPNrQQsiU14wrWqdUPOe9gGFfxX2yldfGqW64Q7Bv5a0
BineQjy57Qre8QqC2YeUN+7GSfaUsV0J1RxIekPWxEn8rPNR16YWfRZnj2uEBgXqwFXevUBdWVDH
as6Z424n0i/8H9/uURMTZdVoCgrgBF/jUBu4a6HCLAW4aBqcVpNNeMMu2kSZL1Rq0apRVFwAyPWL
ped+v6jHU5OgAbV2BgNFp10RYoXQhXd8vTSN7ei7SckUbVZC6pzXJAILi+UVQXRM9T2XpL8N42fq
6e5Lgt43d2iKhaIVgfczIVP2uDdTXJAv3nCnbtLrmsH2kruozX0mD8WXf/T8MkoIC8L4WST/2yd+
jdx6d43nVBjYy9+N6iWo3dd8cVw6FIpvQqfcRPsItl6dCWH+g0gMy4FRBUk677X895Gs1Rd31wEq
sATFWsZ3qDi0bT6X5pn/jDL6PRHhyzagHk0jQcIXt5icMEoMSc7rfVNlzFmiRzDyoMxDwgp3RLCp
SUROMMUhmO9gwEVPNhcEIguF0lnuU2x4qAb5zsghhM+aW1crG9IBmlhdnMoKGhkUsvqU1gp6AkhD
Ws4m6XKAUzKzFjckpLfo2VJLSzvmSQD+vBfEN73qPb6EepERZCt4OCjL7/yrZrVgs+oW1RfK93FV
Fqd9jIvnRdNPKXrP+eeNI7PzZpxZvBDuH/EQl/UivEZ5xWZMjYtNlFw2pPSmrBbhtG0RuVWc433Y
FUaE+ceRjXxPL7Qeu9TzpkxdB8iUTJD0Qdcy2NfnOWW/26pCWA/BaoVdmnQd7N38agGNCvNbMMsv
/oW7WIZgzYTE1I82jwMBR5BO1ukuhgh960E68/uKzPZ0bWiwBg9pUMHm+ak8Kva6gIAWMi4VccyC
Sk6exuyP5LukOJulOKjqk10x+mKIUPzDct7eZyWQEMg/uwiMOI75BX5dOgIoMc6X0Hsp8UDrf3U0
ZmPUUfmke+tPRQBYPM1txHMhcGyH2rlYnOJyeYtp4VYzSzEiFAUaw5smIuvmS3QBCXV+n33U7IZl
fmlrnhOrvU6CcIUTXtm0IaytYCF988axak07f3HFy+eRLvv5zy1Gbm/Ve53IxxScebdy39nUj4UU
HorJGSYupF99+b7pZ7wwBONK3Y/LsDTyIjcQCsfUwspz6lOYrnqY1fDO4izU9kbcNJSmQ0jA7z9p
/in04cmRQCtvp3maGuCA2uLPJ8zjAdm+BnDkcXlxWvolmENu5W0oA4+lqrs2aUplX8SK9pqUl1YD
wR+qMgSq2f7zqQ0smF//YVUxDFYA3tlSjvqxncFG4icFpJcUHPDjL+X1eiOj2LnrBMQA1DnFrEa5
Cj+4rzzLOc21gzqxziTc0WfIAgT8J/Clw+GvGIpLpcl8hrNgBhb28vSkCYzh6lCdIakVJgKIUqDw
cDMF8uJlkpqsj+eidrgix2D4bzNMbGePAfkLCHCt8KITNU+Y2QU324cHjVkSAHDDEIJK5BgySf0P
k8nmHOzmeynAz1cgM3bvmhzsBeyTFnqyLTrVMSpekP1bFLcMXumalan66qvW8QL1jFrhW32DbHOi
IHtoxeRGLBk+wQCIPhN7Uc3ilpMyKKhgGYxgGPKI8e7g0fjbyuLvdht2vzJTRm7X+X556Pa7RDJg
trIITZVBjS+FEw+jcgruBXqX59Rn/+xfHs9w989yrTFDcW10g97neeTfMrBQCX5FadTmGkZyBavX
gc+MiMlNXYa4N73CYH9liJPl73/VfYjO8KuzCTfpgz3YtW8YQJzbs0BjvryrX0QCInpxZkaCnWjA
pqIstZa33EvTmZSCsPDZvZi8C9QxXYQdPlpLIYl4trXoRxi3drgYP9Wq1O/kl6vf9QuuDH+WwSxt
7Q4QSQK9/EeH8SjGqn5o+3QQl4OQWgUsadOgFAdUT9Nw+vah8OT1eSXWb+BclDb8m005C9G6hsw1
LrfM70fv8tHatHGUEnP1/Hl5Ico5z1sL/tpXfwacZUTLhEjIwHrxPtlZSnUJOXD0MU+2KOhJtSeP
z1FYT3nnu7mnF+ymidfmLLDPdnTll7kb/2heFNFMV1oFZ66SaV22T9tX2sKVoEQ6hRXu6kHJILuj
vlI6S4aQLM9zItaRv9CvJagR1oY1y2g4m2ll40l8n6o1vu0PIG/0Jt98khhkRadlBVQTlcZETwFK
WXlUbdQ3nwiqLklmpv6gQs4wBiSbIqZNoHpRJcHj9P5+iDCi/LCSd2LsdqU63qFxKxLqqT87IBH+
GpRtNyraswM9s8QdV0Z63nyEsXIA48dgLyieHYom49FsjbxGUo8sLD55dWAoa7DtEbhHhyOlpurr
LSY5nb+D1QeyYONRDq0IYgtBYF/bckSkmYUFI18XyrtsxRTFs+yZ6yJEe/NjM50wEeDDKcfhCjHv
qeGh5scLjev7nEG/R0Q7wM+JRIH1AONd/73P3pdtUikMMlrxVY4gVymVVqbFVgEALi/mGy2whS4u
HZSKjlxOOKcsbqp/WjYO6G8pc1hWX7AdwU9AdIvOjfzhyRdM5emPOHD38TkYhSaJwCnat6Pp947d
f6RE3p1xN6Iso02W9bfvXms47pH7A0+lRNqWRy4FpstMPw0IHTKFndZkBSfkSzbmE3oOGPFOBnWO
2hTVQIwYVSfdK+1i1zbPIakb2Vk2j7rgVH+486cIaS+29MCIuirs+0/TH+TJCF7Gjmod9cyQEHeX
q9xZrKOIJILjSq6+SK4CEFV32HKDpKRFoIbQUi3WDxMhjeljVRFTNaV60Vj4nUlnB8D2NtwkXwxd
ZupL0GwmzhjAWqKe5XxIBXqZj+5wQSd/jcfH4sJLdwhjy9XldwzrBJoftL2ayjLA+sdVAMbQqf3m
AQp50TyoD8s9lHGM2W8PV8DOIK5APuk7FH+DT+V8NmgJxi7VNZoINayfnrmgQM6XU495CWD4yO4B
vtXXOzjAgqdjQpk6pSrL6snRo13kVS0RKx9X/yeSQvuLDrb6JI7s7P+EQo3PAdQ1p66ynlveb5cH
WoA8+jXUnlQqKdaUE5BGrR82D7Lr/KcTRkj83pXXnPKKPHEH5y0gMtlxDc8ANmyyghtwcCxLqaIb
7lPw0waXFr9IV70Im6cC5UeynfOz9qf36c0+ETMnU44d9zbUxhdelCGKh2MWSM/hAO5ejNQGlPtq
qJNSpe01NzIwZMf+TnsPWGZi7RULei4P4waGqBCR/sUOS975/WnMAaYncnJQ/IBeQjQ/or/SviEv
4fvT3QASD6Rfdt5V+6i3l0SIwlQ6aXD6eopOkByrQBzw2LMELxCyhq/UB97nh9P1BFKzZrMIUFSQ
+pIbnPnbDoCSE2PJClvcPI26F3rHZ5sUEQpdUtI4b/qHM2ID0uL4EQ7ultVa33GoP2FbOHW1lYLs
yGaEVtgGtxyWy9YIT/MJuVpJ1eTo5ECca0NeGCVDBDHxBf9DCDRoE07UcDHnWquUbOhJvgLZMFQ+
qYH8tVGc7X7Vs5RmCO9h+ufJzwiQhxUAlT1uZC0iAHETy2sPXRhlySWpogUHymHhwOmr6Nang2AT
sUYbKlmA2XDLl0hGpbmbBQYJjvBjeb9sgfMyqLOAt/w/M/EvZDzH8rv4qRHRtD0dpLKVMgFlksng
cVCZZV5SE3TZS5lkxjZdKXqynBz1kWSr9Ym1Y2oqeTzXcT/A/mwem8n2NKacPzp+01owNPXwqUL8
K0+H9L0XUd4410kJiTRBBMndb07OYDp9VbM7wdhFEa2SsFo3UdYPJ3VGrehu0l6agk4w4eaJvz68
R6mPCdeXKIRZJArmZCv1Dxq4/dry5iLsglNSsOi8hsIKNWHLKPrSrxT3JcM02MERGSx7bbhWtDWb
REAIi1icIxjbQJsYU04bCo7VIndqORv4UtQDiLDQjLN1GQ9p9GTYXmqe6qBhpFrgKZL5tiGWbeo2
5hPkSDtLzY6Gf6Oeaw2k4wwAliWRxUYqa60J4CUemX8NZ594T5Zjd6gGqzOtHYgmkJ2Pp44K6Tvp
RlBzHJ6fjBfLx8qV8AkYTq/Grmsw4N8AMHTrz+hcVVxZ6epE60HePpxAAKkujXvISvB9wURwAz57
i5/FM06iFiQq0TQ1JdhUYHcWSGZ+MzSuFo7APd/PZo56VDhTTSiCt15ODcgZV51fDtHGw5Fwt6ub
qf1dx6c56ULn2GZkM5aVgGNmRrXVrBKVZqsrlTxpiXF6Kb6n9mX2g+5xCgO0se1UclwgRw1w/Hae
E9MSsJ5pLUwk7/hbrFFlhsGjeBmvXi9VgZVCZlvfeRt3t4rR/xxF3HeypWU9JzocpoOPpMQjufhm
Ldm8pskq3jZBDEqIfOlN8a0YztmmLBBZq7T9kDA61/QU9hjMUQtlS5mOfvzDMuQfrc4DslUJ9OBt
14/2QfsFX91Q0pv0ohLlYUd8HM2PQeB3eLFcjbneVnu/6H8kcuTPhShp4YshFr5Ua2H1JooEcejE
CyExkXMTbl1n7m0SRs80XNybMfedKmm8QdEvNwtYOPFkzg0pQBIvmzS0HVVUlCA2yqxqHdoBxpTr
zRyQQzj7e3sg1JZ2uYSR8caPWVEUMRJTdi60QuTFOmPWVWH9L7okm30OfK7Wom4WpfHZ/s6eOls1
RO8BDQzZJLzh5+ZVGFR2qKqv1VbCVUR+ccOjlwefRASDDkwe8pX/kiMZdUFECq9lVJPU62oTH9Iw
1IdRR45LuwHLN7f9QwVFk2Hb54NtvGr0eyb1TER9/eMpUXYNEPbAR6Wn4HBRoldGvuFOP0teSiKo
nWditaylVb++9Gmf6bnZUTgLB4B5dX1ckvAdyCVIJ/t6CMU4yuKkN3nkz1vtaCFUVNNgumQv7I8T
sThAiJuHQjtnXpB+24q2vDbamVxJvf/vAEARxM9/Ja0erlJ5ZsL1/m/oUHF39fcAuYWwvCYhre7A
15tQMwwLAZIOy0QpLuNz1TTf7bw+1PW83C3+e4p5cemQiikM43bsShftGjb8uxI8dOLULoaQM4MM
U9/qdv3096AtlW1TeZ1TqO9oQZeBcEqAcUH/9n1FrwHn5MAZMkg3nhZD/01Cqrs4efOIuG1I0Y3T
3+lu3XzpxhQY402y4M6xrcGVGn3ew3nUgy9nxlUO+LGJsGBIpQfoqf+kuLaixI3nfueyfJKSEb2h
UAijnBi093Cohy3e7VgSmithIDUv3YCBGveHwuimixvgjhtyO4qj9/7NCmv0kvxLQt31RTC8qrVA
wX71c4oq7xuFbbTkSYc50P7n6VyUDdkWRXgNXJ4N+oRRxApGHQfjXUHqjLOCP4XKLsoxGrFYwftH
z071CGMigx/pp3k77Zb6YycqZ759DdJMn93uNPW2YjDbKjzy4B21AmwaWrKMT0yc467kBvI2Kb9x
LBCPD/lNes6W1szYsJuYjzbw3VaTbuTr8Sf1oqeB4xcMgr3lvMjCNTrAewMm1aziZ79z1PlOpeHE
4ytVMnUbi5rl8HnABPxM0bkzBLOuCF3SbzsWUtukDSjhHKmpIMLtNoG8rtFUgYO1YnqAlvaSTOZr
nWjt3Rpa51+FDwyXZKJ8p0dc6+UUhiCP818Z+WaB4zOFdrkZV2hWWTrB5QJB/5WCzVBVB5JeDm56
UQCL01RVNlR2H6a8yT1JhcJS246LvfW9HZikkCWrfJ6nOhDPO+9GfI+5tT3HX/EhwV0VmhMnExaX
yfoyFQvcwkhqDW2kbIHMa27dtaKb947M2/ggmA0SJb3/LmDlsF3Xh8/9Nbxm4qrIVyiGnGGSgOKP
oJL5ABYIuiAeuRVz1jz7UzL8u20OdcQWtgxKpfSjvEkiNtwn9Pv7lx1ASP7ahsnGKjkmcrXRsg4h
2sEWc4WJpMgGvqeB8oSvNyUuZfQOgGhG4kzS8WawXu9rw6W/oQftOcEEw2N0IylCoq57RUVuXJDj
RHkw/ZSSlaZ/DB5cwGX4FzYhrtwPapd0ab5DjED71M6cy2QfmgJPIG0cYJpO+ycEKl4loGtaFovh
YVwCN3VXAGGJGUiOkQ7REHlwbKzTnr9GWXfKI0IBz01WYMp7uG+knenT9sb9uXHeaHiGxphlm3+r
bcT8Dh6sY0ppnQo84xM3V40xyaXIqiQBPKOBO23LZ8S4bCEADRN+Otd/mHAoDb8xTKggg72VFlkA
cBl9nXY8UwmJesZYhg2z3CU+Pj3TelavUFH6uScmvcOsrySjaeUyYuUfLRQcnvEm37rcY3N/IfDP
13tpwyEEUs6rclPBGw0Pcp6G/Ra51ocDOBljJYuD/GphjbgWBwOJeUIs5ow2cIY9q2ko4osXoJng
bBao3ZNlu7U8UHyhBxXF0eac80ndDy2YaxyZYdm07/0cfjNl+vIfqasmASJrWSh+jFSabuuVik8o
a+Xo2bWJzepDxXihoWKDF3Kk4WYuszvHi8A/c7GhrOu9CvKcwg55/3C5wtMcyaX/wkXPF8ORJr0u
9FCxLLDdoCCNEDO4cKHxLaxjV1Igc84YXrSRH0zFEBcxg7zoTfr50nOozYgPlpeWZ/OCGgxxC7RN
bVPt8yjDJS2W6bIRTtWE9zsNdlgyMmtUhBxFARLLNrahebMK0XscJPlbkQTOOdWbrwHqmr6Rozcl
2zBhJB+je7IaJKCiP1Q8WjAcrt8fQMQuQgTPqQAsfSusT7J9e4prcN6xfQn5isL5E8sjoSP4+FBV
uaxtNkbPgNXJQzc0kWapPrRWtcA/7sk6Eck6K6viv903Jvx2gQO684od63+uArhAs66Rq9tJd0VR
A5lOmcrG+2KG7i7zRK7yqjo3UR33ERLeqRAnXTwpqwbxRf5OctKG+gBH/a7wy9v9rhQsZgke0vuy
ry5AtZXFgZyldFBa3KLmQPXTy7J4NAzgOJnqWGQRlnEGJb5OulWpR1JHawkig2JlC+gD3qDMuYBs
W6F/sDapoQNrctTwXOcudy1mFXLbho3KzkcgusndezT/AZwaSI31HsUADUECAQaoihdo7bc8wwym
ASP47FJkHUopVsI6aT9Y3Lt5914j6H0keTTb9UURaQMzgNMEFR7aMCrtDcKBAhhnISQrnDSLHN1K
iTLkuaTXpiZ3wk4wE0Iz3givZXzrJ4dDe3wozZ2g3HUGqe2p2ZGKu8/2h3Mrw9Z4tKgnS9TiW+C2
fk2AYHhDyW42FsIW8EWb/SlaDmjGATd4eJAfMlGWFFaOAfRFo8av2JsbdjcG1+P4cinqIebOY97v
vMF1Dcn4uq3Yj2BtCLWFY6l01OgCFsAc0PYerF1tQBiN3M+5rylMFMvnpVAeXdNA9sp6OIzC+PWX
vBzWmlItbFChXSCilCaOQhgYta809sUGELYVJksbdyzRD53ndURcGyzEWSIa/TBaVpGDLMLP7qYw
fCgBIm9LtPT/EDx90Sovh5dU8PnfG4azabS+/TM5MMLrV7oKXRiuxGL36BDm+75VEI6H7u+MkWeP
5y5ynsRVgmywB9Z5wn4E66qqqIHSzVOGiPFNdWiDQuzSIFKL7/NX0zXP7GMzUKjxoIZGFqg0+AVJ
nD47ZDl340J/kOtxJVeawCHl1WubKWY9BQJRYs4XpeiZy4/w/6mMKyrWG5JbyjDQi2bXa7RkHC6+
pNioJKeeP+6FpmLSiJOZ4HrpUlagrR5n9oRO4DxHp6zSSzqFKO67Drig/G2E+3jYANUQHTYahdFj
JUrt8B5iTT4pWMzThIpOJjVYFTfmx/r91PTheH7IiRltJO1avGaJDn0QndCJ1fwuDLFwicHZuxPq
nevNH9KPu9V8LPTLZQZWXMbad827xwZ82J8jbkujZdubLkP0c+l3CC4R/njCAOIgSjoL/DWs9/sw
6KuvdY8n9DZBxAiu7SztrRNk5oLfrfAly8bn5japCruSHd55cMzXb0i8gayJDm2UiqVTxSquRQPP
MqdbpE3d5BvPLDiAQlxu+fbSbX3M03yi+ut5LWR+lnhE+F9ojt7XyiLz+qHCGErvVPnE846UazYA
1N2dGNKRYoJ1MipnbsTZEcc3SiCdoQJ6JIXJCGvFO7odPssA26zo5wR54hOSuMeJOqmN1wB9pMmf
rEb+wev2+Mp9+NiHNIyudJB90VAptHS9nvaeoCLaZX3XxmiznwfNvtbnr5UZmnGLgQagqoXeMfVf
ZuUimVNhpECH/0DremgvU3ubwzB4dF6yB1aEwIuJUp3zfPt+x6nkU+sSHGEzvaFoP3G3c2BQrd6x
YUMniLt79klJRLQNO6TIICul1d9P6KmrkwVVZItAAf+rcM7x55WkV4B2Z3eOFf7OKaywykXIBvA3
SBfD93MSA6FdaE2z/rFhu7q/KhSFSEN1dnnhnO687u1hGzxlBMW6mLQo3fEQB9jpnyCtc1hy+Fvx
GpXLBs4Yc6YobEw++Gk5to/D5jZpOPongWYR5ZaFUQsYh/A1RSk8Pml1MhJ0ucnwBxhCaT7CNL+A
SGoixeJKI1++IkumX3DY/zMUaxST6Redk49A58kkSRQrVWhE/h17xklsnJkNO6EZziYU8Tnwmdw/
KJYE4EWGcxQmms3tEKgRx2WwgMY52i7d9rYh6ocMhvIfVGFGwh524ZlLDzkKdc6hWanzK2FwauY6
/7okcEMZPGcJbD+/oJSmqaaKtUtoEK+NwQT76MVhnv/GVmdhcUnBmovQgCN033t2BPBhUxRB6ziS
F84Vegu74xFbc2+EL8+ogCJHX8Aqg77EFsK2x0M/ivssCnn4ZGZh5H4Tn+UohjyY97D0/YV8Z4KG
6CQ/u74q7i0w4+glp1EWPOf/+q+02/uVuBd/Zg7q2FYyJ3e0OSv+Nrq0SHFKVqMwhQZc0g1YcbT2
9USwTvwqsZ4p6uunakA/Fnklbq+Be3l7IOVAY/D27CGyE82ikYII4v98rN4X3HDDNX7FPZzypFOf
nDd/zEb2UA4v4BXEWTbIk/tjC0UUseDYvET6/36bUhWQoy/rO7Rq2Hoe3tR2//4PunwLS+tuQd0z
Kt+swgxLNk3enYTjjVn9mle1uV9yvmBh9+8UE4nxBvmz70OQ2amwuuARLaGrcqV5JZN1t/ntAEcp
uyOyKt5nz8hCw71h0z3pS5XemsUIKuDtPWsJZu86zCexCLrArUzcgcMHbShEUPY2fXpuyj8tYRd3
L9tE0PfBpxRlzfS5cM9EEuqs+PcxfKKqJ+TI0WWTxZ/9aTyuhA5Grf2j/sKxV00k/yEqZpko0NXg
3aW/Qd/zoW3zQ3HBoUYMQk3XEBK9XYlfNgiP8po/zekK4PcHCcWS/1EvBol9rb89U3LEPBBCS3UY
ACRTuIONeUl6I7/Tm+dvYWUep+RhmeikD53hJFsBZ2X3m8tgHQ3J7nVij3jashJ2Qx4LeYMWtfoj
7NcBGAzufkFpRowlwI7RY1o/V9GmgfQePwzwKdCaY/xfJ+8219GkipwThHStdqLh5FdVsVDlfxUm
BWdAH4ZmV33dTH7XDmgWX3aqnBRozGeV03qA2ZudLZkTmfCUAUe/TKoR/aNhO+g2Xb1L+xBcqdjQ
I9K3v3Swy72mk3UQI+LQjff4zCA62Ef+e5WTXXAV88o2Ce2yJ3+oYdNH1Ts4/jcSGvRqYMaVK5iR
1vVstZ8JmY1oxfaY2Y/6vBdD00LKvsfWdROXMZY2tPK0gugJPEIeAwoV0GN7a1+dx2gUX6A72/Uf
WXQ60bIjYSULc87Yb9OoBftVVg0sNwGSeVFEDX686UU5W+wZDaDQitblI62uv7Pf5cELOMfmwdUN
axBkT7GXj2jdpiB+DGITRvm37R7fppvmAF/EMtlURIGodZc9g06vQtxKHXnyBbybOVLxT59m6N33
xXw20g5YQDgABJqx82JvzkXDPU936VhOll8N/z+5XwxSVdCFDMFsaEBpANfpzL+eVEH3HZosJntU
BAPQ/hB4ApqBKws83QmIbA8lYhTIcrZzlxjAgOGJtcLpCqZIoUjpWpFWSMdnGc+woTFz/est37NI
iB9+HofK8REIRpq0Ah631YrEQ5+viFZQ3PA8CM0XomiwZ7/JOPQ1GbHbj3mfipusu0hwqj5/KdzN
MEJ4jgBAu0lyGfStJtau6bVf1Ev6ucTC3Wh0V2gDW3nJLYh8GOadvcQGeHb0R0fE2FcY51Y9F0rA
1l07I+7WhgDmbBCIzhBBADa6LaaN4dh4wiIn+GDCbLC4aDZ+rkOTP6CdXle816w41AJeXxDVhlTK
nD0thPTuC1AT7qTS6QTGLWls+dvX6c7JhnozkD1hjbxqQWU7JgujsxHZjPt/Mli0FpbNC9Cpqmuo
q4MmVgN3fHAxAOTISHtCjTY/Q0AxgwD2wljICavKaWdEoiOgNxp0XPB+MNNNrZSZAbOxo9oVf2x6
YbbQQ4FjK+d5D0FVQ/qMPfZWALcZJ1JeUZDfkaSKX64VOV7MfoVtlzq8HQOV8uWv0851tfnfFUVB
bs2shxxVQfX2ZIYoBpXohjpohOtI8/adCzifR3/EXuFag/7Kg6DnHaxOqN9m2HzIMbfSBcZA3ebk
8vrV11Wj8pH4HX5rRtqTJSZgq1CtBM+nA3Bi3dQb6TerjDRfSXsvOQYfEJFO8DIjK/p+44c2dh3h
3/JDT9fn4JxuGclGcvsuQT4vJqyQQ3C2vtaJVwnob53IXtRIgky9kD3TP1ZqilA1Ago+I6fFTZqW
LLYh0ZTz6JrAgcQ9Vik1KefyYXfnP7hj3u15KIVZNik1S6O8m4onjD5dqmpQ7MzJ69Yp018WESJX
N41NA/5+Tv0Ue52AeljuWcd6cD1IUQPNw4pQWG1FeDdtrlw5yr2o2B1TDfbH5t0KQHRkzLicu3fq
Zwfwffl/O/E9n/3yQ+wZaubhuLZQ1z4MUKaTcYDN3Zgm0DDfnhRTtudqYetA+WvL3wReW0oIvLvs
nImpq5shUOx4me+N6o8zvUeXBrlV3lyS/ZBuDyiKeBR7FtJfh5W3Bfbf7JmYYFZkgjJRo/to+iBB
kMRfbPe0/f1VK0Lzfnb57aNh4pfKZkRDqdoexctrjZIVLewiG7KrlYBDHocSKPCTdfBm9DTnZtQL
OGcwT14eG010xpLFuYi3soB/VGsAPfc8W3X6F9cSA/NQzxn7AdG5JmTfNhYOqZxsBdj2ZmTbYM5t
34GlDFiGTijGE4zW9a6eqQ5cS6UfMw/hc19gyH8DWA+BQ08NFsYeBCW6Wb7HU4hzIM8VB/wGnH9O
yODcC6TVZH/WoF+9H1Zvj5kjF2VAm3i2mGPlNof1jBtsAxCDEHuwOIX7F1YeTrGyCdPsLp740a0n
nlfCcX//ryQdbAFfdFxpJkmnTqq4qkXE/28mYeUig5e48VKL4uXbijm6r8+X/J74ErqvRjdkRWOo
k4kiDI9O1X4rwqnVUT3xdyPRI7I5Fph2SGdeisNZh21O3zEtjNHJ4mxZWqfJYoJEZyLnAyOkmCVl
2oPl4pMY3BHk3WYZlV41NzvQmLcKn2A1CXG9nddbvmNDCmHky6uGdG5MFyxFjL3lKT3Q1rjUEhM8
mtcBRQPVe95IrgBOyjTXOgnkcLICK5Rt20LwBOFY2uNY+rDMV7GAJp6C8W25rgcj105gYmdG3q/7
cNrTfFUjdRmaLNRh+yR18Khr4lvEzXkXgkedMkgAw8nrX6wwnPoDzHmjOrkqjs/1ZgiH4yY+xZMb
On7P4+r6CSLZ5MPU0gFkjxfgckc3BUXLXpoLNIe7lTu0mr4ZOhlxTg7nNnhZxkc4R8NcYmyUAIcT
BEgAc7ouHIxUJt3nEmXrnmOvAUyUFV/3Fz7wfOg7KehdOQwhaMUuyXsFId24dafF1Xrn5fPuqqUf
eQnLTwjBgdMS9IQRNDUALh3x68iEhXrvEyCAthIz5o0mDkemG91FZV6sO6sQV4+JPclYgtVFOnnK
gRqoMEwYATCEi2HjEYEso9H0wqsxgFnpNaFFQpGn4lFG20zc1h7FHpc0qtxQz7wwSLzwGx6WuZQW
/hwue1VHvr5JV9h8B7Lp7xU6mDgOo9vDXih8nGCBz+Ppsnk9PpZdJ8nj7Uqb/NfQxzgHDM7B3ypi
7mbC1uDwP/a5fIdz3Zgcnrg+nNFVkUOIk8psS1rGAjR68g0fMErPLP3R2/fdGkEGyowP+t3/6m9P
UZi1Yaji8EPmoW/e2rMel1GC4Nj8UcU7SLWnwdic+6QO5AdjJbkSOIWPxSPUBBrHY1RkPrvyiNP1
21wo/U9IejpEEWcgMRXrhRDfO2GpC6IzZ0Rn9879dr8DUAUvJWiu0V1ct3CcGqMIvvVXust62/Y8
H22svqOkC4WBxfRDN/6MtQ2p8rPewvJLfKelLTBjkzWTCcy+EDDj54OwLDmpNKLsbL54h0l0ktwL
d0j7zX0NpwIC5Xwxfu6ffo/SIYPyD3IrxyRvpPDGnf1zHr1mubNEOarZSqkNm5VbX01Y30ypfWhI
WSSC79Y4AEYsSzhJK4c3/ZOTN53zOsk4F7qWn6g+mPxbWrk/lLtTDbJJaVQrJIjH4WK4A4CA2ZCx
noJ4ndoklEOtfvnEy58uytYCcYfl4Yabj9FW86Wsi7d/DfZ2tRGRFyaUEdRUZ9lGhYlLKLF/FE7K
tupEVrCpBXjjWK5C6P9e24xxFHLWiEJevLMI65VAosWNwTDTpj4OxPWEQt7YtJNcX9LSlWY4tyu5
O7Tuz/WcvZpFztk3lORTNuXcdE7k942C5/KK2hGliJVyqS8eAcdZrOMT8YvUVrpi5bEp8usMpCRk
jHcCssHPw+wqFILOk9+bHpuWjUOgyN4334VpgFn2FzYHknICvcA5LqSkY+fb4kyfo+RXZKpERE8k
VVpeuwkMHxYIoqJYIaSp6uC3DMV+OKMf63vOFwAfJvTXxQsdvgIUgFhpmnOrHfui6NlE96XuQX8K
UG0bnb7MiBi38vIL2muleX1xTnhobBUA5fkiCqEV4G8xZ+EDnnz06VLB6AYcvhXgJpRug9//qPpn
nTDZ6F1Nfx5VuSYig136QsEewgjUOLxEb6kD9/4W0GAYqok3cZUMDZFJeqkRq5BvXJji820tiwV8
LwHlkFxdPFhhoGg23PsILAgBTophocN0yxpnJgZkt7r99eUlpCsYAcaUG0+BAA31BDg8vPNDKDnG
aYMf/uuyvS1zcBATTxEB5hYgmNeaQLs70J73dvgBeQqnHOF2EZWqbEVEQvwTWKjhtpdxAuBDa5Cb
FjfM/sQq4Hhn3ceVTpFf3Bpt490vLtNkCOMEplFeL+jdZrbSvvjnFetBfBZkeKf3VifiZyBTRWr+
pxn8ldSXAclQvcCwLhQRL1YRVVmkeACcnQ8ueAy1p9bE2FLqFAwwG51/1SQ2wwE4BM5HHik4/JdR
OXej5NAqb52PMHj99dZVSVyUO5874Z+Enol3jMpKPtCJAbUkpEqSbd0JCwvWq3xF03b9T3BIQL3v
Uo/1etsw2l+jnN15gzvxuDoOwfQHQnpxMrFrIb5CkupXsQes3EFj1Eqyme6o8w8DqXcrdgiR1oYd
/7XWiitt19DkGwCd5PELlXB2VQKG0WH3NOaznJUbNHUKiKQr43idzQUCwM3nM2kBaH4whBCgjsPU
czEmeXYamaZS+PmxTsWhZmGZeE3Y/WtoOoAqJw+h5EGeWWcHZxsGpNrL+5AOQVv2juVI2zFv+pqa
5J/qiEiUAG7nLkwDGugA33Us2ARaOsthqnFPLcMlWJx2iF0A9WX8MLMPYT9OaC2jXqL3/GmsU8u3
B3cNj9jhwPWP5I0AD0nImgKL5RPZNF3GDUWEjUI1yfllJD42meqlQjE6rVUedmvwu8VspLs6P3dp
J/YesyzN07eaoHC9zCA5S2rWORkmEbmDcXU9YK5L3nSdN0mCVQxJtIhmbwecoMhht0D5DZdR8oFQ
zLptkW2uk0nRU6OQuIsiuI0olEllVVNYwrq51r4cwhOZJr+RCkQRKfhr0xT/GeYbtHOeiIE3sd66
f65t+hprWqdLEhpBLNRqye5g5B6OoGukCRupber86ryJWDELVzGxg1YmwY/DNHNq3gLMt6ULcUZj
AkmGMUVgmLkDl6knBdu8KtYcBQ9mRptMNCSkZ54UYwH33tPdKVFFak8YCY/h5VqN1U5TcJoaqscA
oRohvZHtFiGMh6OjMROIZk2f6wN3BrrAfMNf4z7co2dSDVk2Id9yVj+k7/BElF9Obx7rexaZQVJZ
Wpk48WLEt2t8+vU2ne2bu+es9sv/KvFArBUc0I/yTfxCruE1HJrNQjJ7YtPpSlw3IlLloT+Nn8DN
Jjp7rmsAjS2dPk/k39TY/Em1KiwhHVkEZSqK1P98QNZ2l8P9nMDOgyBgaRr77hE9kuBCr6WTh3jL
TniqkQ9mB62VvauByijO9CfO8ihX71/nE4upt4SjY4ssbZtq8QuhqiZHXb1UG3VvXn3zBA+sVnQ8
g+uyeQX8lkXhhgAxW2Q4K91vrl2GOM5cEwjyHHRDgqsFTgJ2lLrqSjaT2Oz8sOfRUJeI5TOXHEnm
yJU7RYLIYu+1GfkSiYmmdU0DkS/OnnAbqMR9xF8AsGbWDCeg+PXFYbU8WsF8QAQVSmcmPA6t+BQC
MMIQe9bJNjW+n/AlN40AeWcJVn33ThAvQnzA18+viVNusFDYKv0BUhVPatQH6FGHM+FqqPVX3eri
xJHkdcOuNWQ8ZFQ0cb6jPHIMwcDgupAv/IT926qMUBiOwRGg3Hu3MRg6I88a425zrX2K/8uuq1BV
3vR7FHdAcnmjI5ogSDIbWbhDj/UTO3DIrSB8+1z1T8zDq4iS+yFhXHv3pDP9IsSniPKo3YI4mQT3
MwookLWNGZLrK25kni3deEBV3uaqGmoiSjOD9FZzjNctZTQqpTstfjV4Fd/Uj66hQE6OAp6P9DCe
Vtzky/3iHLyzIKz8Nl95ip0r8nH4S/7tMk5JbHVgbDDjIHntb/pgr+fmeNcnTOqy7B8CPcSi2f/a
ubzLmytdjrDO+kLhhTLlp9x+1JU/2dCL7VwH3em8UZlNFgE2mJQLWBcRVZ7EYPKLncb6w0Bi4zuJ
oon9TNa9EdRSK2IGaK9d4x44xdMZxC1wAKzLFwsGHZ/EL3EVyhXtaq4FKFLHWsvQNkd1BdMKJ2GM
P/yglWD2XJW/Gy1j+6nJW1f/YC+xnQqrdma/OsKY7w2M1wPTuWgUJ2WFuDoTUWhjOZNzFeWMbHa5
irXboWacTjnKT2BU7SjrRIYu5GjPbW28xuunFVmL6RWxhy1Q7WYK3Ivhl5A77uG0uwc3qC+yqmpS
ME8QG3foBcK4oeIBS96kB+sshs2V0KKCWE7he34GmSgPBRQyn7f8s3Ht+cQeQossP7aAH5Dj3Dx8
N/MsuaPsVho5Zhf8ZgAgMMKzca6vc+oT652vYiOZg6PdQpPhdjZ5iK3tG+FHaXbRDX1go74KT9bT
5blc6QarHWtonIcoqwcHkcCNqPRhUpcnFRsXs1sGUQMbl0iSvoX5KorO8jO//qAggeuC//y1qAlL
oZXeXKFUjCd15Agru5+QEZI/BeMeytQ/s7yWDJRseWY2P2S8Ecb+Hv0sGxPa3qi3gr/vtXkPmrip
eNA6blGQjFyOaRQ0brGWQ3LNUyRkFY1w7tJsSX8AU8Jk/5cTsPl+arep12cN2gp2HuNcKsVA0DJY
xEL51dBmhAbNnae6IvNSxT85T7148OW5pacVowGoW4fw7IgzFCH5I0Sh3oaGFX71dVeluSPA1wzo
gm6NUE2wurSn9upvqtzefwSen5BWB5tU/SSYW2rNq/wVgc7D6y6ejcB4Xsc8IM00wsvvjccYBZ2p
Foa9qD0iau71cAFP9bBFPfwrRxTVTHRjB+P9RqrdwP9GzCfySqvH0XvHGboCx85y6tubhNsUu4rb
FH1Qi+0oetjHmP1+Vl6laKyTyhGfeBChoFGK6qoNBRrS+vjxWfC67C6g5081G7wsquQ4zl/xxWmN
zgZvBp3RZpoQ4WoXVDRnGykXC4gjSWfT20IKWFn/LVkKkM+vpwtOlP0/ikDKeOvlDwesD3j48Swm
oImZYjq6u7mMSSVyGdUr3293I9vA9wurewuhuURDbklSkY+JCyJN+0zLifLRWaBSG76vWSvHyv3b
JA4/gjepACOKYYPCmZniqVacndcpq1WyxPiv9GA3ERtPtFNqaFfsf4Atqiq5XaqvvWpLiD8RX5gQ
LPa/DZDSEU0AIKKreHfEs08hqO1ffXHOl960ScPmp3hsoGEPTe+XagiJV74FDqetxnlJVI7z4OXB
uIyep/3eLGdcHX5b7WWCjDTQRcdCcK2JnE85BAXcexEHXqullNevQ1HUQl79G1vplkziGEomoSn0
3sOFK/CQ5LS8Jm5cjcf33nuNAH/s9pt2dP2bsxvbHLyDyyuLveMvYdZrFYsI9AmiW4ydxWG5fpTA
2/hdGkRGLwVXOaA/IWO1AhHha/dJt+XdLCnMgSZbVARTeDZZDbFvBDvTHnru9490HJPQS/9b8Q0o
7mudk0Pv+SE2iU6XT25RQ9GuMGoetT3xtiKwTmNRP7ygp00oJL4y4ke5Zms0IzbsLHQyVyiwAwj/
Qft9xamwJTNIKTlyhLBcpPlyjK6k3yNUDADrMRCgyQdVh/mwFjlFbQ60Qr6bzF6fUnke7KmKd8ib
WPIoFkUQvF9kN96ticmktC5ku7/qXEyOay9zo35Bc8VALqOXtaOlyZnQpBpCIJPC3FOOi++PAXbG
G3OuNuBtvDQQiRKPwV9DbBKhgptunR4cIxae1kc5a62YcCJSz9p/rmmDTnztG694GcSHMaCrtyGx
+vfpVb0uLkXswK1a9gtDFtfCndfnlKFO6PXB0iV4zYk/WDubkMXMK21iQOpHx5tRXm3hv9hbuLD8
lRoZ3MicXTwKPBwa2SwVRuH5NkiicH+k6jBJBsH1X0LQvttMWl6II6lcYM7QH3LAfqBnxYkKhYKn
aRWdZvfkzLXiNxghXa+myoumMHVclJVVnXEsuE2hlTVlkvKnG89jfg8n8ZLP0Sa96K/SlALcqXb2
Z//wAz/Uzr3DUWoh0hZR7narzMEQsBgYUcR1RVqaSv57fSoDYzRLK23Ol985ids/bxzuEJo3GHsn
dXTIpl8Ta08aFWGj3K8KXbObbWssjad11OFDGx602c3lcZBSumoUBSxPvqqhrg+ov9/NskPaYgA3
8Yp+8XVM+JNkg4JcaFczLnO4DgGCqDNDaF+yBofJuPx48RE8d6sQhtMV3vOTG2fBQCXhlw2JPN1y
SiBpzyvtdC7CdZGDsDnKAiWe8WV7sgGUA3M5ryBoji0hP78fSzTEjWaJQXcuVtJGMOEwojIA9KiB
bAcXUk3Uzz8xMJgw98o6RXJeJCiG14ra1ZqJhO0fEbUBX/Qh1fDXZQC798ocJYb4ALyD0OKQcw9p
gaBv22lUvZ4NLQy9bDhZt7EELYPTvVAPrVazAY+QiypJYZWJ2A76YaKrBsYmx+6q0UrqtTi9gsv0
aKID6JRNUV0cDndSsltOZ80duMRL03esPPTehPEEYsOdWWcgCtqwiL74Dchal/1pgMTFOHH3q4fa
9AcvaTC+PqR46itYPJ4D1fG3WGwgz9xUEpkWHWQ8rtbRyjZS9Y6WJeWy8Ecav8R79fXC4npcgDzU
XVFAvQkkcM97jmPt4Q6xxKkxK8hrp901lfkvPWXIVwX4KOBZXZaVddieTkN3DukODb0O3CA3Gs9g
ZRJykXXBIEURMiRbEkwVHUGz1U7Q9Nc6M4XKIvCEns2mEQqr8FvWs3xb8WaqD4oLqWsiac8oKxPi
2gC79nYaMRgQWkepT8W+2peMMCjOfKUt8mpnvWPSveiOaVAIEx//ziNR4Re9RPiVzl+DfaBcleSW
/aNe5aTjgnr1WeLNtVksTHDcAqKa+aTd+oZ5OUPdFPJ/qKMC/mp71s1g/RjOM/XdmwqrGW6VsEdo
GLW2W+fYw07ZFUtl2MVxX3hUFsqiZsJKtGu63/SNHpsWC8yAZqDUcZSBL2ppqVP88q+2NvRuFnAB
6wiQ9cP8duP+zGWfXYWnTJ9VC9DB1ZDAgPHrxRqlEx+owuLp/zOmakFpHITCBnlhA+xDhLSW4stu
7zuBWYpyBJoDhBhsywv2NWlKLeoj75Gu/KqL7O2pGhQ4LFrleafZkc3q/Q4Q5ZY11bIwdHj1/LJs
oVU2g2/sJQRO5QrFOK432mjyCFiqm2IaoFvgmVVOtDjsxb5PR450LricRqLiatmsFzZRN84zdMgV
IEHu+wgaB/wzyp3PRS86BofL+NiQOCbOlH0+D4sRGS3vKnfssLK3FmUbsVx2spx3HV76uFbhpmtz
S7Qej+GVCSump619ghA3HYWWrRHx3D11gAYupWG27xLts6g8Gpzx4WG6CsyQyaxF58REHr8B5K5G
xENFtGv14Vhop6FOq8X4oD6zRGwrnh3ABCj7HXuTt/uqjVKkuMlfBzkN2/1gf54qj9if4JUaHhTK
dnWK6mclTJ+qtE+pvY8gjmHINW0k9ouSQm/4dnb75lhw89kLMO/HtovcdMVG41ow8G8OVBBT1ZLu
TN9eCjcEISPk9QRHYphQiC7Ol3Yq8DmBCXIbzP4lkJk9bP+R4DNa0MmzPtM9MJLmdYZdptzck/4K
4dFhtlZ3HzvFIJLEmf3K70x2OIGQJNdnEuh78dnjjK7T3kX3SS1JpvFB5c5nZvhpwHH9/d7KwZ7B
MqnFjen7fx+kT4OkE1b29c5Sfo7ZdhhdWGTH2dWFkkCmmLcuyAE9Go14NSmz1vPnSwscBFXBvkLv
FFQLGCdTFwZ8NZx3dgYTlRv5BOfqvuMp6PAbMPZjLllynhcKlfbQakUn+sHKzXew+Cvv+70+dUx0
aDhXvt/MRJtr7gysGl6mWhGPXi692Ev5snFW+7L028JeIyiZKW16EYbCmXacBGknyxOIM6kknNMM
eanxZu9CQKkx9x8LmT/+IPySG8zBMug0QLYTuVs5KB1HTWmuPND1bLms3BGe4SZ9dL/6LdoUJSi+
H5htWuqf/nq+4QF4rBPRGEdow3+3oFFedez3OU/nhzdxQMH4UVnjXkhVBszObu+5cxaVhH+rIpAp
le629Swh8XU9IklqR12hyarkhYorO/gC6demJfNudbFMN1AqA0dOC1przrpAhNH/U4ZE15a0hlz6
ijPw10bOfhFCJ1Z001K/aMaZkOCvPFUxcyzNDZJjz4xMQyEtP0CSaGIRRTF4mQwNBM3wilXw6TH7
BaJOI2GRCCWNyn5n0IAMJC3dSDJ4z4CDfergtHQty+XlUcPGZc8LZiwd6onsf/GJER/SlsOugFzw
D9izoeFH4XHGWO/F1/j4tUvKAytgJAYuFAuLTiFbBqNdK6yE+1CAdnnxO/FnjubiVhzVQZ5NTpLZ
G/W4nt58trTP72JwaGP6ial3jerGPjnMMyD/CJSEmQtrm1cSnTkdnd7RXOxgytHVUjipF5IOCVrd
WJn7/pa9j7MVRsZtgDQCsVnUqTl4y39LHH4HuHBJdbNNKHVGu8EX6nSUQdbIelsnbwx7LseTirwC
OBIeJMM6HFOB4TPHvMPNzrUtqGn5bwuKaWo4asssG0W/uvqBGmfWo+AJdns/4sL572JO4HarXj7K
f3pE0l3F19NBa/M4iuL6BU9xonvv/66R1KNbzEoSGTI2HCsCumsDCYLgJOGQX4R3Q0B8x3RXbS0G
aWI5c/7Fjf/oS8wewPLq72P7Uh978BM09MUyr/gMnRKWIhNuFNRr5uWcRc/BpV5Vp79p/Smv0VIA
TPxYHyRnc+Wt790u+GhEkVACGDsfdCttXLvLK7ZD645P2QVSyXD2vL8BRgM1jP6ejs4lygJczPUr
yXCC6ig+VBImud4igbfkiSIUk8Z0YT/YSVbz7g7CrWHNHotBdb8KFA2OqxTYLWdGJSPJKd7bhHE5
96bcSmC8csFIHqaXQxf1yEurYLRuY+ffk+u/zzS891gFluIVW9EytwrgDpfmlNyT4DhM8fkhqDpR
zzFc20FJlkJsgxzeIOyJT5mBMRfSPzkDwfieeMTuSpJZkfZVPixRQbHioLPmDzO3lK327gHhSy7V
gzPQ2rU11B3W+D9kQ1LSkiBXFDXJlJXZlw3xW9hvB3ubxQ14Ya5TW0TvWZqKCCa72bNsWIZbml+U
vANO9BAy8lrl6V2RzKZJjHRiq5j3YVKPPIbrgsOrK0lMvDrpoOfnjgkRdRPzs41eE+nRk40Ntu1Q
pckNpWxPlTeU9lgaIeNqcQoFSdg8ObHQDSBxwH6+U0jO+gAJKOCZYoaQTbyoy/YmcDoZAqhXr/65
fnfU1vm7Evs1hXpinVBR3+p8C7r47VyEN5xyUX28aFw7mJbwhH+ChzOpYrYq5JLkPPvUt8WIcM78
sIdvaSfCMkEv25+X/6fZP7N4P/LtVayBq1HQoEwEebDUWCm4UAik9gGUM/e47VEOiwBXKjPnG2LQ
WjBmM6iYSjGm8dFqEdsFUhs8/Qz6/sKWvZCNoX8FkHNsrJ8VBGGl2396bBL3OsHOU/PDujtT2biI
1ibgvYjxesZERi3VgZZ5bEhajlwPAV7/ajL01liuUYYr3KlPtm29aFjnzmCHKMap343bF7uETtJI
G1kughFbFfuKFaJGKvwKV9ioNzcpWMsjGGOay9bJzd/VKswxAgrPITnisjk+/MVqPZU0JsJgVXpe
cL3ibi90r0D8/hHZZXX33zjUXdeHQ9ZsMkyaxLjLoLS0fJO/XlgSKjRh3o58rTeyxOPOD1QyRKn0
yNg9v8KwIXcpkgxXU+F4c9CXWM0tNxDsOOL/X9z+X/9xs60+oE0dQqldYseywAdE1SFP/Z4f1IzB
yWdRTgHVPz3H53+JewSLcPNcB4RXq1LTCEXqEyBHAqGIagcycAZBh4FG0jpHh2ropz9cO1eqqcC6
95iRMaJW1I+50kfdD4ZNtkOchp8d68B7WxUl7T7uPh/v2Xv/9wyRN1/8O4Whel3i7joY5dT/q+25
sr2x2nlMwIHqCWUPI2rntdBdHjUO0OBtipAqwrpmsxjhXSe3hxFytGNlXqWch3MDM55As/Ve3EWI
Z026vlP+8rlQNLbAmsQDDCcPeW40N7SkaskDyFrXPAJ8cObdGSj4I+7Ms3ORh/sP/cNM99odHX46
3QMYQwqZP/H376j3sAbjMib1eXEJbjgqHbRqP5aiwTe3ztY2z4hjqXmjiUEU68/kWh1DODUqAoxf
LA8hWQHuHPtkpRJClPicun4g6qH8fNUyBGXwHa3G1PE//Fb1NCFXCxAlsEIE4gfJN+RitLE7OJnw
y4fRlBa7stkU8Uupxc0ZW0cIv02u1vRc6nhW+azgZIQ1IBgE4We6+HvM3DUYSj8a9P1TwMJsFTZE
6+uZ8jBdsyhah+gfamZbeBJMqMiEGluJATaKCbqrsvAWjdzquQjsAmD4CQmf3a9/tnw8q/bo+Otj
sr4/5/y8+XwOVZOZ0Iu5MAcfdCBwGlVQkbCulF/P+7qQ1zMNU1/uZBdGIHfW/8XmD7s38uIpdcHy
tnPA0bCUAFBBo/4SwWNkgwDYMrfvovTUIa1Bsgbdtpe6z+HG2H7kgtna0SES9pPS9c9EuG/ms02f
3n4OIfLKMCKYMC3jbaphLm4btE7R210rdCOpSU/PTrlx0ZMwxBsNoL8IkFyafROyjPb+tZ68m31Z
/141gqmfWJzwSQxxBzMa3+ESrVY19tz1NOElde+4EbjhMe6bXK5tuouvABvp0QA0KFvIvg5cuEOq
sn46N86C03jCXiKMhsbHK/9M4Y4TVV+5Vi5TcgjqXpde2aFcS/E/bbrr+PP/713BSaS1uSSuCjGp
DarXqM9exBv1bB6B2FAEbAl1ez8ZoGYK8iuwS7RSM6/vlFpvqRqTxcMD6TEklMZqlXpBvC9oFU/X
SZNfGnKoClz2I98QLS9u2O9CgGh88Zt/p79k2tAcvX1qSl/e+U4x8quKn/2aqIdsk6RZV+9KJJx0
58sPrXcbiA4I2uUVIzjCH2eHFhyJwIUJMhDvXknmw0JeHytrwUweKOqlk1qICzTjVRImrvV+C4sM
SuNzU/XgRYZeUoZuzT2i5k1lA/KXlr71oVSM/oHgVRTxOLE9bsgMvD96n5OlPWv8emAPcaa/o3wm
imYJcQTVPEOufSVIH0jEORttn+gfY+uWbPvErVZfm5cpl4CVZRV5wzHP5CdpOfudGCQ6A9cSbWqf
0I/gkL2lUEWP0nMFUvPLfY5gu2si/tPfPl18jmVosc2rOQ16zmdKXL5YJaHw5QD1tYNMBNjZsrYi
9tapDBkB41N6ZITxXfqrqPzpT1yItVSNcgZPARRX1efsHCDJGg7vm21KM/JKGlro3DSvqhHalEwS
Dg0clogqL07AKMJYEAaYD1Uo+1PfNuMaEbLiB9px5zcEkfCR3Oht0OeB+Kkfj7ThqP2xVQ7H4fB1
TPrltLxnzj6fQbyxBcf8HQ5SE5x31nQ8LZD3HttsvGM3fl6mtQVAcPdJnWYxlWQgwblxz3XR4F2w
uScmzdcEHH8hO/rfk7ivCfdbwY1g++JBm5kBVJiLRjXadPKL47i+Q8gWd2nQA2+dE/ySF3pmfR8B
mtzbjDAKAKMEawGsKyfo++6derCJQ51mJW/DYjiST6HZltu1V/9yyyxbLJoNAfl6MXZt01mP+MB1
Q2+/tF9TdFy8ZY7ZhKnBFE9yByrj5ZUzkxXNVKHThpnMUOPzu9VWNrA04gHlMFvIwNdmTyBQIJcv
LToWWmBLRgInt1gCpTRA87/3N1vud4LA1F/qksptqXEh5phV/tZULIrgtvv16quOEa4m/TMdKxwF
HRenr028XpxccMtVS9lsF3q/ro42EYumkOkM1Hwh5juBjIFtg8RlUpc8PJ/blcXP5WGyEkjmXpHd
lUiqvt8ITYXLxrihW6Og5g5YWv3QRBVtsZ3vGLYxShHaCqCjcNC1bDVwbtzLjQeP80kPO72MF7Tu
ORDvw9PFtlkWYav+JTLdoVjwGeLVVE6hxW/8HHSr93a/u5kZO6rrk18F10FDHqr1qYrqVZfiNnH+
KGtlJ4LZBW3aAlqmBabOcZ9bXq8HZuPFId+//x8s1wTzdX7rXIVhgQqM4/W/c/G5SEZXHQMYiKS6
QdkthBNkKajyX3Rbt2BITfpJ5o6HvVS7Jwfa2ZSOI8qJrwPV0qvdvUXx5wSoiYuYXMjtEoEyEQot
bMQyPx0jyWDTpsCH5Ov2jMe2IyRjlbnhNJgix/qvltlaW4O7JMUc51ROcA2zxgrPByheoWLFkE5r
giVD5ypkNotOkBtplUTfv6V6nGCelpN+zC9QPOirlTTR3Osi9bT++LHLL35n9/QBw2K0xr0Kb3s0
05VOKe+Po7dGN1S+uC/c2/lnAR3/LH+wCtsgImolfJ7FowaeOjutduz3jEOJbMvjDLJXs86lq4A5
Ow1gtPcOykZrEw1tx9U0Z8oBg2FtVO+tBqQOS9NFgVijs1A4CRtTV5XEWzbKKgOFHxeKuC79cN/i
xfoFCSTr+EfMsTxqN7b2nH1RldsZInODgxvv00xITg8YgUKPhSp5Xayb9c4LP2YqIpwCpTw6noOR
hO29YOmaI1M1F+F2JO9VZYsUU3vw7OC4TUtLcK1yOU2N3VlmJyGdLvU57Ueol1y251mUox9KWgP4
XP3Ai7v5DsHSN02pPcD4Hmo9ThAJW3rAVjoSG7+93FarURFccKyap5TTRJzMesL2Al8R3DY7OxeM
6E2MVmK9+Ura7LCMOyPvqdrqYIYBrZX/cEBM1xhEdwx1AjS61suiyqx9LgsYBunlKfYiuDhu24Pv
4mkWR3aKkhM+jWCRWPhpaJu0y+AB9P2lEj9J6dHqk/7Hz/Wl0LJ5dP/u3x7SYFp64Ebr1SjkpEQE
7eL3oCixC82mPcTv3L88ikxK3ynEm7iCKa/+5JfmbB3VI897DALGevuBBGR7cXdurckbl4en5HGV
x2qKLQmDT2cq3rdSu/37RUq6+Eu+zUI2+y9FYeJJwPDyEv5tKTrp6P0Z/2OK0ceeIwiv7dSRXUt1
dXa9rUwf1nS32eK7QYYXWL5kXsw1OonRyTdksKQxL+tgpoh69UiqJGUoE1S1csVOIPeyEAwELPEc
wBNyPoVic/Z4gSF/mKSjNkl8gF9zs0MsCi4M+rVFaZwBTUTAQ8aTF1hquYSpSA8QnEGsL/t/cA+h
jmshYeAVsh69Wgk8J82BVxBC4N08m/hwBi2twfBvEAwkC1xtS25Ne8uVUSizBMV2QzGD9MZ/K0W/
CajIcVRykjyoxQot7EQPLYeCaG6mVPp1aERAFIPSlhHF6+7NbbAQtyojJ6OPwH6/0nq5Rp7T/e/u
06BDEAxdhEwU5cg+0VX3JWc2pgN07Uuo7SVHTHLhHiF7Wf4xuMI9xqLqYU3CO3hPr1capp7r9v5d
PgaMsPRoHseCVj3Z3gSqV2+TJCpK+s0AyJqY73I4rI9GwEGlrJgkslg1h1VRA6XtPM20kJjgLFpg
TAysJadK+9JVrK0PvEI2uSE1tNP5nAmcNELIAfzpBMvOQ13MiC/gIYNhpHeEcd9odDWo9va8DVwh
SJcCnehPcoEHUADfrxjVfdv0HeUAcbZbskIEgjKGGKn5TrkNd6qVpy3RGxTTfp0H/IAaRoSqp/YW
q3UvBlTWCLd7XVL954Dq7+UcIkyMkeVuvrSU82mL6KqdbEvoXi/z1bPko24Sm8h2jgmgJglYG5PP
HUYjvX4JyJzLKHepbOkVGMbP30GiTdfmrQz72eiUbp7n42pjwa8P5X6epUqipOSgNEF85a9NJGGU
t5M5rm8nxcaXqde/vkD823D8YOKPd/SCYK8fehTq+PtElDYHC7tFpk6lrKuIGotFr9ZzjwyP5fj6
P4ipT2I0NzNA16nCKwyyVW50X/tatHhS4QZaKdznqVDMpLDqf7DXBSVmyddgdOwwqe0i7gjY78+d
n4FwetzCPrXyobPs+1BRtmFCLJH04PAmobeSrJbjoshjnS8PhuBKN4/R0ewmHZ5V2cCgZ2jPl/Kf
A8uBNPqE43cgDuAvI6uQWuL3L/JqSTjftXdkgZT0DWRpYiaQXBvcxqyOjBHT8M+PbmMpxShPHwpL
N48rEAG4NWlA3n2NJcoU47EIc1FX+owQxVh4sft+wRJBwh73IgPjmRCgfRURQdF6Oz+nZaKZgtxG
lLStyqK+DuHT27OimAXoJ8ons37mqUAcLOiqjCexDEVvNJ8GwAx8IbfS/Z8yeCbaEtsu97rqOkGg
AqK8LhWA9dwxePEJOykS7K6zXerfWuIl+QdnaGsuKgdpiDzd3e0QuP26gkDWJnbaVD+6z5E30jbm
APO6sCBjbzh+dqCYsOqDUIgIoJvW7uAzmSU/CzQQIydUQgv+z++1Fo3hnIwPn2S+GMo5bJrbhc/Z
zr4WIVdCap0dyloD7lDjsZlLZVCy9gHJ8XgkCJetqosSWOIRY5aJ2En6gtiYuK/m2njv8OEArdF6
vWU8fvKUlUlhR2I/Qr1997uxSlTqG+Y2FhpYKT5ljPd/xNNak3A3vpzMS/7iD9im0xD7q7bRjT4+
y5R618QCQKmp52dQJbmMtaNl+cBHxfkYT889Cm0ExYNcw1RslNH+NH/IfZL+E3YILBhTiafyn0C3
GkMMEyBGKQ8vXwDevUTnEoPeWV9FHwF3D81OKL7XKJXWUpd2HOw/P6nicQNsogBo5TYeHvXaZLZa
owoUG/24Vs5qqCD43df8qiGUYALzZaWzyE6KRsUzI8NUrwDCAO5BEmRTb4lSYh9PV7DQRoSGh50+
zs+hiR/9jOT1YARBSuiqWCx76KPH3oAlH8vMxOQTVX9AT3GSeWIZpzN8egoeQrSrP9dIpbPW+mOv
m8MqgNEIhSDFjOJn2EMtxEuZTB44zvicy0rg7kHu0kWuUoVOoRxKupeXduzq45i1daHHMRK9v8I+
956SMXp0HAFVDt/WKSF9P7uHsMe4yY0FDCbbJpvjgPtxYPcdcy1JNm01cCbNAWB6n9dV4cN1TSkp
Dn9KfsET6eWbrEG3OTfMUe12kFFjfrvRXGgofvQe5OXxKi1/GchNhGOEGHiK2iQOGRD1HQ96JkI3
EuuGKiy17ln+MyZGq3PbzQzNFxfH1YjRE+RV9exsHf9AcSqmm3TdBWNVxKUKYBiCpnslX96q48zY
vaJWTcqajt/i03YmdFGCJz0zCaeUqNbVsvIy0eyGcre2mt0B7+OzFlevl0ujZ6nTTiIam8meYZY3
TM73/kaH9GTOKMyKLV9AabW86Nilvy+PseVEm91c4nOxdyYe/Yf655X8QIk7UlX0DYNBv5uReZnt
N6fuZXsuq/fAPydAVuthJXMt+HI1wV0vhBfE63t3ZPmTsFZ1RK7UzKVS1oQqze8vd0zh7SjMeiEN
6IsjD+o92T9e26GnUVRC53lG9v6m/d9KOsozMap4hrSGUF1KReSdc19I7+qYip9yZBXDkOzEqRw/
hfEoRqGtnV0LWpUdvyvMB3Wa+Dw/h48MVGBBFvHuINiNHAIq2ztbRXJTKNR2ykm6g1ndACqsSPhi
jEeteDaxBEqC5xvtSeq8a0ea+sBi5wWTiObAiyxMkbrB2IReCrOVefS/oxK+R+fcGQFDAC/4o9s8
UEjDtvw76l4UZ8ULz5/gSC54DlXa0qt/PZzFkTCGrW0dm3hk+RrVmszkmzwnMisMqJXnt61EQsdR
av5OD+09NCG08r55VDetJ43sRGLooe3K/arqBeTVFSKapaY2qkgdspOn8A8iZhEV98EwVzZiZXLK
UOzvzbtsBTD49qys8MYtodqfN4zQu9N8p6hUmM3SMDY4y4ycmofuUGHMH2x27RG5sELBUu8PJeJL
rmYmlur4lncnaHE2n8e7u01aXSjCc18O3tj9yOpGQhrvgDR0mG544xDazY0NFmDLo3Uv6jrIbxst
Dn/52asLw05ODfLmkeVasddjkCOWvI5NT01ugi3tTOUaY5eIIgwoxQDd2GKhz+ebEWUgPq/qyyNf
dVtNIdY9IlI2EDTwGO+s/7z2bdISi4Dmj0G6wVjpQ2K6O4wrd20BfaRud88UxSb1vNa+zpahWwEh
o+3/o87EzeWC2mG7Pty2BfgKXdEv/BTTZdwCoSlHwb5yYADGrn7SSWUiRuNlN+qs/LmArht+a+c7
1irFZK/n7lmigwzPNkRG42x0vYfY0UOXyVja05eWK0GAXyGn1rdtjVmeLIPatLtMblIEtK3N7a2K
ua4HXa3Aulu8utHmWWwff6OWsABtpaVbUkEKhti7BSuxyqDRrOt5ipxjEbIw5tYhXKlv/YUyhnVT
5OUfkQ3W4F8bOM5843Kp20gjGE5BuBzKsNYwm808pnBwUVNI9HPSM5xNlx0qSg/4gDWAu20htZfZ
qI7BwZseDwL9vsbKLTbPDXd01Gw3F6FGnWcCgRwqL5sPZ/vL7wcSCLncgy+XyZvtIpqCm+SYgxxU
lFkWyZLeJkp1qfOE5D+eNBPbKZhkrvkmU3tfO1oB3ARLYsYkxWN+KO/F5JQ3VkPTi8RJJuy5+PdN
YRldBg73wWo1vRuOpYG7+Lb7Efa2W9Qc9grGny5ud5mvLvmZmmToI4XDHn0zgtWffXTZ6qCB4q0O
ntsWHhDeXxSFJWJdoTcKEShtbbwq8JfrHMd7dCEkGtYsMoekWwN+YDo84EkUUee2MLwLk+GevzCc
Ikcltivhc8F7MYq9YJCWZeGV5844Nizg0TXsxgQ0gKOlpYXKv2YVs+XSFc6byM0bCXpWz6d3KQhb
nJdaSRd5QLqavznUdQSuRX7V0tn0YfrPotSmAxdFlVt1+RM9ZGbz4hc0nGyYLL6yl74tlNlzPcw6
bdNeDefOHXnLdqgsccBWTOoVC36jOKFU6bLZhdQPZfqjyIrJ4Vp6hOA6xb1ItheqZ1Vf3Wt87ia9
p8kmHUmeMNMSeXvykwJtC4XboradY9ZSMFsxnm5cHdkE7aVVvza1bUTvieQuWf8hJbBtFh6Zqa5b
BZVhyQEvzz11R+FI6yM8Uz5a02CrP7KdDMo1UkalxWbjaLMVPpWjpDGdKCZPLk2euc9/E6EtA3HG
JNZCGt1w2/mdY3t15bpyjnAL3y5CQX0hvWL9K95FPBpzx/ooYRmTIny5yM31J88gnmoMQFvyPVEA
NB8XSTCUtbVefKjd2j1OuwrCANE1vueh9f4E3krh1VuSIn3ZLW4R9xUDk7F+3WtV3Qcq/8G6Zwh9
SGZpwYQSI/K9WGTcifc1cBCd1MH9Bfuoykgo5M1yK1k7YZVX1zHrf4IPLDct0Pzzw6j5b9wL37Gh
+2BnPnPeeOoBDPEDCkfRpimqo4FIrGH9a3t0dGFKGyN1jdcFJxtpVJtX43DojNyiemFSuxPvqREI
RZRR+RfKC8USJ85p7edPyPBHTNH1afkny1EESWsgdwoLKW/lBjoBL4fM9JHiPSJL0s5XM/zHwbWa
BocSNWY0JV56ldMXnnEpF06eUYhom14Ee8CyuC+zTsMMZ6EEMMsJQhryq+rv2iL3wp0bFfwaH3K/
wXcKsZWWytb27c8E2/1pPouNx2ci1CEiiPEzb/fL47jXADPtQ58Qx5qImq3DgB7Ssp9Ec+t54Ukd
HrCVOSfMrCKPp7HWp3Jq3OEamDthnd77PSwq7sffI+rXVP8O2WN6ehuvlvS6sgpBs8yDFllpaB1V
klAXFtvu/wImhertklAkEjKIfK/lqlylO2TndwUtBI23U9lCCOyiD64qdy/3LWuNCq3vFE2H2sln
q0oFEXy/Y5NsinAfwM7uyYfVVcEeKIKXHGm2Ad0GTWmpfm7ApVMBxgW3yUPn3hTHQutN6X625Lzv
gQ6zUPGLHWV/cw3ifBH+zeUGdffMiJAta4Ca9cVS+ISdD5TFfboQSbJbZWds7s9PMbLfPyPMHLtQ
YgjtAO3f54L3hEdJ6qbZZmW8sLpdEkcGwr1yzygp1TQ7fMi0lLKkFKEnArSjuGYSN1aUWfGSz4Bw
Oc3nxnOVCn/ja6cJoQJPJmIWbWCAW2mABEKJmRUbWXaX4jKGPFtduQZuGes8vXXVmFAyIseVtWG+
p9pH6sH2CnNDjpQiZjsXEVqcy35Tab2l/UH8dfRUkD1HEpIT+gfYXHaCo/UBedHtiv7Xh8SrVjAi
0VhxqWp63FWob3XQ+irG8A7pyJWStT8ZVG/eJoAAzNtR6g3Mcp4LZ72bSc5Mfql6XUBmFiAQ++p0
lOuX5e8Zi4I++/uNp04mbooIH/f/gH/fqljc8XOTaTHbLke3lV52RJwyk0UhRwjSU3Nr8JnhLVZn
icGFy24aVw4XA6aNYCMOfXvgl3BqMUg+wD+3LC4cbfQIyNJddSjvQK8WWnJgGIY2gTa+qh2xhUB4
Q2akOufFrrnNk8CE86FtLhHzVmqCyK5xndlSPOocdAcsklQCIKCAC/U4J1bTkRQlulAcBxjHtCpm
KmGQ6kFxpvJS/ya2U7xgz35AVV5CovtsRbqwJuz5VKlFUGAH1K9qVpCHnuh/icMdhCbq88ELts1j
FnPvajR6iU+XNOPFwwE1VT1rflzclyDvYfy4QjAMaXauW8K/ZZWkLsNaPe/sbQ0SuuHekAacmLUr
FLWPUTu8Vne33zw1y3RggJlo3lCmOX3UlYy1gIaRTgorSzO8rp16VpqjvSIilZMxWje+3rmlhHSM
xcSazPaanCDDZwFXlKbpPDZ+GspnKheh9tDOo3sy8fX++3QEjWD5EsKTYQAW80t9F7on+OiYPP7k
uYSYOozw8Ll58H/2zrmFWsvShfyq5Qvpf76S1jyqK/rEOx6LR71mrVe8/QEQXOwjX9iM2qP/gnOI
86G7oSd9Y4qShhaLLdGfU4GnE4wxe0PbqVYyKOfusTtfeiByF9LGNZBWqZraoJPeCy9hxo/5qGiE
e6/fmEEVIMTWbJOfg5fxYJkbwmz7maAcC0/xpVDiIpaIF1wyS/PMahk6SEXJbVjLlkUyVxfnPl+p
rUI52EQtxsCE3vDk1nJm+6vWhXVyLbJf1lO/K7Z4B+fy/oUwBpbNnhzX1XnL/VyakC0wSVgwiWM5
EAVvW85DPU/odMNwdNVOhUNznCjcdM70UHPSlBsVib3FiCCuNCOKbNUL8tofTs1cVw/nqtwPllJz
77Jv3AOjs+KJQqYSN7GKCEKi7vce++NMQj/eQX72BsBS/ZsRmUqpdiujawVu5z/5K3hkcWVEaPj4
152IZyhDYVMdeoxxwHUcwBA1JxTRd38j+WUIYgxsCZSUUrU5tsxBlyImvRI2JFyI3v13vFwdgGGr
X+WjZt+jfnif+d+bcn6G+IrgDMcuRAjQ636tTHARNKjGduWCOVVhA7v/9xPe6Z5xZv9SsOSQ8PDG
o5QFCg2ELLwQn0Y9S9t05MNEqmgRHWDSLHiFsbwaNJxXyu9cmM0YrPO8r63PyT9cySJA3JVmodj1
s82bEckAR3hYcb1Rn07N0vM2cGJP1PcXwuXTK68Xt7E2NP99hwCQ88LNGbGgXVcp/7rGT1GSzUmd
59Lg3CYyuDkEOB4SEER5DhPeKzoc+2+iwjtNtln47+mj2DPDQJafR5ICqdUS3LS+s46kkG3bNmoo
Zww+02qCvGzpJHLb991zksg1qJH1hayLgdJdBQDlnEUFYx4+TWXb0VPHbTBvmrMEZCxbtSFD6SlV
kAZcNjTH++Uon3iRK2GFC0JB95f5yPJ2OwMmrqGHE2Mxwxj7gh3YxIoq8CcSBMMaJR/kCDQTyHvK
fKC0CA4GwHCZLiP2z1045NC+pWAFak9OhGtofN3KRUEsPEfZTyeAfY8wEGBLv7eMZvdbv81wkT1U
M/T8qkvzcuIGqTHFYYgXb87/nMPNZZ5njl94LJvQx6Ow316SCEvHYlytP2HDxaWwrvq9HoQRawnf
/Qm56zPp8OHkOn9Um7rmbI/2CXpYaHJcCExVA6D63/cQ+YYUSnX3yNg8zWAx2QF7YQHHfA5WQPBn
nEojabd4yxXsWUDKBPw7K3hcZ79qEpSC8YXQO2oY8tpERDvBkTeJGxaA6a8FbjWF3j+9+7fgB95+
JZ1MZYT7u2Stx6AZoYs9nyR+xJCxpMOPIhYtyPQqbMP7vfOCiZoHO/keIPyI/p4yysmwU3CUsfyO
lCEyVGtgeIetYs5GE0xTFQ0v+b+dzxgLnl8CFriZkgi0hvbAYftukL+SRiM88vMinrfpqzOCh3sw
SD0AusiZWpxay470PBtwDpqKWeMQyfXblezK6oQxDFJnn4w5e2w+nb+1Zjj+XxnHv/iNoF8HDuzS
JVh1qZUstKalm5C8pkmvjfm+Wiccbn/4zW/83yFsT5k4flmYRsdUcc0fkfx0QcpPR7mLWymZ7p/j
GG4st4aNrzjcX4OVwrlbSoSqAiqPQStHA0ohxtsKQItK75/8nMmAOMyzQ+187EFc96D7Yd+f+Pmu
gf2MTJMTKurQu+RnNcxFzIN9AJoItKA7KnUlhbCEOuzzGPvV+fRUOCfzxXsh5QomP874SKLNjJSV
fbCBTm/Y2vRAm4Uzaoo2WSI9IHDXuKe0TxOjLDb9eqecsIykLujpzq8pFJwE2tILLFktvj132XR+
CVnioC2ItxG0jQxrOIpyuNcKUBz5vGyPJZo4U7n4NNwWwMMsM0GIqQ2VR2SXxDY6DG0JJZFSD4qu
PqCxq67Z6wr2ly5jks3dgo51KBRktTmWEJbweoAdpWVY2XaRVlEQ2qVp3/K0Rrn5F/4UUjZd9lfF
AVfBj7o3HNG+7j9Z8NVmhZMJKqaTF5NDWWIWyJUBuhcNkMHcsjniBIdlnPvPBtFZ2nPiOUSA0h0y
+zWcZDnMEWDEeRv/3fRASkdPwUuZcP86qr3l7QmdJQ5MP2sd25T+nSBcAFk6gSguGNzsTEESaGom
/T43EcXl1opWcAOT6nQ/5b/IHOOKWpCWkK86TIkBk2nzlb55cC/RqGo4DBXP4POkux+fenY6y0o3
hz9/o8t8c48CgTsNxyJupo4l0LQpbNRDavXePORly6O0RRqe0TFMCgxPDVbcBJ3AAeFrJEB37UBr
faYsLsEiuMd5EuTzmz6B/bjFcuRjSvCMMJY0bqQljei+buYw27bMp5DdfBWm1VumZr05wBT/1kyB
tW/JnvmTN6LN0QCn67M6Gp/Xz7OiSwZk0fOywAE06sDdF/RILxnA3XOYjFpfE4SA/4eyd5I6xlTQ
RPhQy2alXdxeQkaDfsWLU23QmpN+A906SR3N35mSLG572y8snhQ2Mf9+cpSaJzWAOtHGul29esBW
8lt5J6gVwkCMrzvrbdTlx2sG8IABmwdgBHmFVdJ4te3OMMxGoHxYqoK5NLdAte8dxVltaGPvsW5X
WWOgN98Zn48jvRNpN0PAzfZIGC00SIO+pzp7icm9tO6pSH+GsSzLHZchGWQAaAZbV7E0WkZt53KN
YSCefF9Vq6WbVIF2qqbglTocZRJk/d5Fi0x/JqSglK4TqmPMcXo9m+3L2w+wRsEnWDFGMK2mjAki
0itte3BqdDoOKVsuO7POhkqZrDgDVDYQNW+fovGN+2RcYEYy8bAGG9N4TWt1AWHzxlb3N524+DbY
VpTnIlRjq3oKSdaJiRuCQ3+GHIxQ9iCYE92DBGZh0aXjQFLYqggXWKWrova4p0i5gpaLNImkcM6m
NNV28uKRrxr6O8EqvZpq3PCjDt//cJzd7ZgzTJWzUGPH6fhnKTiXFvc3iQBC2aOmGg5f/b1csE7R
yYC35FHIcYz3gzXm8AHARI+Q+CeqllgHIqNmd2atNFzpjC3mB3XZROVyYnHHGNs6JxvBrkQY33n5
cPqkfWbVikaOw0yBp7n2tnvi8ESzh3wNAcN3C5KoHuK1MB8frGHAhTtMTpglT5o5ABy7/Cvsb6rZ
wc5zxl8wgc6ScLO0xZkT0yDOt9mhFVTd8AYYXXczsb9HwP06djPctca5Wb5IVO0ce8SgddR1mxXA
QPSeBbgUAKEdrbjF5ST8EJjvOzFI+jY+cgaA5c2X2C7lT8fnUncRMOz56Ogp1IBXbzEwZFbKUHO8
/op5wpnNzWMLFXq2vixAklSExiFxoh0b1Mi9SXF0s6f/ZFd5eGwiowPYqdUxWWAS22lC/9PSVPGL
HGmO3+2OsRtkMOYSrO6DCc/1YGbzMiV2180kBm0u24QXyBbS9VbHec7ediXSjMwNhV1YVMIwRMt5
+zfw1n8xoTKh7JO9Wldu/tNYY0kRRQbh5EReZhwo3A4lxF2nuoPbwX200sY8Jx4wTBHv4OfuvbEX
/Kf1p2f3m9KaGiGAGxfyqCMXUz5da9WxGoPVLHp9JKJCZZ2Ra71BZxtY3mvhuliBSYiAatVv1lTt
VR3+kdjs6itnwG8CrarjkpX+iTql49exDHuGgiQhoU+U5h6N9YOi8WYZMiJzRka7c+TzgWrs6ZKX
xALZbaXN27fsDFPg+jeAVZ1j9T1m6+5ocgqKLWXGubcVoa0+R47NQnCw1QUUp/gLth4aBDlLUKYP
xIYFhsuu16LRidfh0knMtxi6P8HL+PZV5GYVLaUyzOWcSxLeGk9MGoZ1svHbJs76QyVPNxu/r6zf
BMSwuA7eDx4zuSLrgbK+N+IjoIS9CZAUTQVfxNt12YQwyRGMvOyFimyGyWv2f4prhxUpYkS9zNXg
tVu7nadS0M4vebaTcKVoZJD/PGUiNdhNrnZC8zBxaq5VO0T8pqiC0YWHip5HYbt52deMTR4QRv0m
ED5jxT61EQGjUdZrVuUvq+w8KCub7qvFg0MUPSrSW6lgPKFmRlBvYdWdBf1GOMvtQ3Om8z+xjO3P
rmwnroGMwPNoR8xZSPD+AMsXQmh+7VwyAkb4vhXCuZZMGDCD00ZinHy+dQYJ+zDI7fXbvTA+DKmN
gzLHaJc84v5iRye9aguSTrQeJdBIxBNGWiQ/P0C/kJOkUS/ys+PDs42bUgo/ATaT5yAZBZRR45qT
PLzT+nmArCY2fWLZ4yNnCxDmJXuogVvAR8mMx9RCtqNj8rGRg9emEulaZkD3aWu0+g/qVvSDS66d
evF/HWsATWyLa3Up/SwKxGEXXq6Y00wTXZdlo/w1DMfku9kVoJTYkDLeog7IpiC/7wvT8uu2YyzO
20MQbBE9fdu+da4+SOfDPxbM75azYhJ4GVjjhT3ObEB80Ds6McR+M+xA3x2l7jx0DRB2sgZUXwMt
r4S4QPFEzyeDcXanmsjoaFBlLmkWn+BQ9KhNuxMVtKAAFEoPsrlHgZ92C1xB8faAeO402yOd4ZOc
91aVMCE7T1ExJ2JUZZwt5MGBpXCsCiIVT7XN9C27rmrjFCFfzVs2UIE2CJJpa+QrHMy6iVmtsO8X
vfcZtGAXT5iThHkdTm5ARCI5ixXJZJdFInxaEdMatORvKwsQApwHiX2aMX3pCCHKxeCe8CUmbdjI
bLUmMa9YZSiAQ+eck3Ft3gCwwJZvjGTK56OP6lBCskGrdplONEbFAc3RvgNDnbaPlN1EIZWdNdpH
6fCdFyG+42UQGuPv7kVWup6i2wDUEud9u12L1d6mYU6y1yDNrwqFmyFffNn+di+dx3NLj0fIZoO0
vr/QUrW7qcNCzQgUFRB1Ml2fwBpRo9hSvX/uSWO0MIFwyUoTrJjKJhtrgxFcyV2+rwB73CCvBcnx
TRj8bTyJ01T8pZSYYojoRhA9UGFNiQyops31C6+5sxsqiiLNhQV1cJF+iVXtFHs3vuHan4A8qt1K
f3MNf4HqNUBxOYgCcO3gU/xAaY+2NyDX6OMOpaXyOHeqgK8mouayZV3XNxAkZJIs78S26oAHuG2N
yQXG3EYxSlOnzfUVL1ZzMnh51msaQc1sJ1Ry4aFDsr8uNDcmj3Vuu0X+2RpSh86zwiGi3N1p77h+
B2yhv5z/vkPwI87kU1DuYbFTQm14E6HS5mu+OtVrgPdItEZr/xwAyi+jhK5i3l8iKG8rxoTuXF1e
oz5A6b4ZLoKqg2yxDqsgzVCLTGRvhJfFcxIQB1sa0pCspCfaAMOxwj0YJmC7U4qUt7Fj9d2SXwUl
QKcQX/f5h6HRV595Qd5SnQ514dhfBiYd3+IYfz7YUU5pH5XIimRwEAVjVsy7gRrk24vAqwcMpmq3
zNQMu1+HHRSm13VChQ3x8knX9WBNK4kPqmgK9smh04zhfZDGHfU+4VPrBLlo1AAjSiobeeq8i23T
ziXU9qdP2cYMDPjCQg56YmdzGAAnZhzT35N/R54MaIaUtfLw6JU2EYkIJQI+tHsxnEs4HmZ2woPh
ijm2qCcrUE8a1pzA60BMOc9tKNyk8eVWle5o70ZmslTSuqWm9zw+IGvBTOhMbmiGwLn/v6YBtlGF
Zsx3UZqq0J8T+cbgckD9EK6EmMwZm9iIXG9Kt6LCw7iMoinT4iP6vaWdZHgwzSz98zxgzN9I3ZiM
xSlTpI3ewd0TuZKP/z1x2hvXSVDV83o1lpEmlHzK5P7zI+uimHtvTfGd1TPEtfU4sjAyFpGVuodS
WbDIDcK0mpo8Cdq3i2QOEQQJcdXbdm4rurW0HyiDjDRmPgsw34LZTrmxzKDKsT8DtE5rbGHOm/Oc
xmnnuexZp8oAMF8JfiYRXKw7Yw/GAvrsmZLxxKo1ZZwvcnUFNMN36t+2My1colWv+r7pdiMi4Qgo
rPcWkv/zlvxGQRVtK5W9qgyXgbo+FlTmqWHwpas9dOaCOl3JVZAbeXWKUq3ZU2bK5295+JgcLQSc
Dt+vWpczMpK3KNwb39mDaeFGxsvEUArNfMdopCVOuSTlv8LtwWTYSEpDQCionZqrzGhvB/i7quK8
/lDyVd12wt4TE1HWr4yBOXYiEi7gdAWThsDNx0WkN1IYzrIO7h7djwPra1TMJGT7RKQRgC5fWHPL
zhjZi2npVrgNwM2wVoskb5XrfbYj/MLGwQQSCEN9qx28RFlkBLrLHVAQazBST6ic6xadLTwhYaLl
efwGh5pZDoC4F/HSY9noyPnqiZcJ2BWbE6L2SRV5T3J3jsf4K2HyUS5lL3JtjL4w68JCUGHN1lMJ
e0VHAgPQthZpL4ITONCEiuRJrhYtkYrvCk4mQzoXXfTgXA4klNCDqz8CPQ+jNAAxuhpf3d0R+M5o
RqO2xPN1crhrj6hf/43rm1yllYRyGO8F8A4SxKuNGScR9soEY95uDXkNXDDEWdW4V08lRJWvkAzf
QoTBRYqBCcO7hlWFWwXnkQuO4bTwDjOt6IplMLTtjG7PkBlCXsqEWxsB1wJkSaE6I94qBCEYuOtw
BTZLMXaCALL898Sxa69RXkrCOM+hFE+4dOnqsPcoxjeWsIhdLkTHSUild+aKqrxReJSTFQHD9TRU
YdHGAKE2Dmu4fpsU6xmi9MyKxnbpsrYkmLmNmg1pL0B2ycBf1OxRWEGppgZ0by0gAudgu+qkKCDf
qw4IjVh3E+SwmdScdjoDADWGppjsokIEitW/uOLZagxDEQwn/ZoD0JsNMRpbki8EvjB3sVda3NjX
m+jRcKlCAGSI5miz4909KHPL8u7XLCkARSE6/LRML68s1DbrhFzwXSO3Gy+oWFxLWW20FUk2zc18
cpVsmjWHGZZYQMsjMrP204/wGY97ky2Zls7JNuPh8o2QX4eDxju1Y6T5znWmnKzVfbQMlKlFBgZI
Ju+jRQypb9X5qc/84/OWMQ6Q5abrhQRiHKxcBSNlrJMguiEfajl57TLo6Pw+u/xbs6HizGknR4wa
mpX+UgQ46kFw0LQkw9FbGIy0mr0KWm8gJGJbYbu3V4nGBIEpHyphR146cB5k8JWh41tUUuUYE6b4
T7ixDzmEWZyUWut4mJIg7gIP3y4JwozP8Ajq9XdX2hq1mdYdbjgJD8TO3Cpd1hQ0jWxj2aPhhJ3C
EjKeFU9EQOEI9xOnKXpV6Xfe4+DXjNh3bs5rv6uIyKu4EI6SugL3+u8RuM62wXSXqxpzRH364FiX
d9dku49XGNjAkhkIOfQky6qJB8E7sERk4hgbs/z/DdR68R3ty+07Rk35eQ/XDh9DVDuvNcLVJWJH
S7ivFoyaKmH9HdX5RbMfshFzunI1kgYE+ebmnS16vb2Q9VicdQVZ+CsKs+DkvYC8QIyC1NCa1/5j
9CE93OHng7+S0MaItw9/Eb9CmUP3CeY9juKImO46G6oB2Ke6nOn7p4iau67Dh0QKjFZPbf927CqI
V3pw6r1j8Um6pdLFo+8mFSiRpEdQNye7LEaNdD7rW/+1mKQBzQQRu6MXYptBIFY2YHyLgWIDogGD
xKM4ZtXZnRHVySqnG3WB1NMQJZyciHPKpE8wLdl9pMu4yD8ZN72H58PwvU3phYej7qU6JB0eaG82
5hmslvlGVA1l65yecL66S4nJGTpnNqR5wf48gD7Ty1tcjoxMhv4xqw3892rOqTGN4FyTKAHgYbil
G1MZTfdolEEHCfnvADQooqJoh8B9nL2RVbiWTmsB38yAUBnjYQvhJTIicirF/gXEoAjorPafsShL
fYcJmAimPdG7NthBA4MySKM+eK9qBeZQoj80Af6HxbIgLr8nWYewNQsZzERHBaYNQjQZ+RdRLGFd
bAQu5cEOHlIsbXCj/M++SV33SdAYbG6BTQfpSejHbnzHTgljhpXvIICEi+UTEffCkhUWg7aR6ruE
wqFFOO2MZLKtPyd6HtKBL5R0Sz40q6Hob8q3mPbBSLMnqXBGocZtR5Al7JylA7ioz/sxAi1KQM2k
2j6LmIo+4t1zCH+MdHyaE4dz9QcoRRiVHnwUTDNRqaXsxaxdi6pd5mUETMFv1OJKSfv1hQ8gLrFi
w4IvQ8SGgWBv06QZCVDTMsU7NIVb2OzwCELiG59/kssVApnAsgY4pKfZkK7KSGV+GvOWQSXbok8g
WTFmOCVIWnZ5xGM+huF7xzYGLI8sMO/tkNq4OUNgTR5Co4+jC7l5X67cjw8i7PtDoZ39XScCUskG
R/LekY1drK1mMoaXAPL6yZxmA1X+cO7yE3RIvUC2V518evqhnSL42qJ8M8rLpYhLaX7JDH0H0WUm
EaIZDnbPpuA0rcQgfNUSvDeKV27tV83MPey2g5seO0yHN2OG/4RS5mKgmpZx6L4yMZIAJJXtz4Yw
9Wct4wI6yO8ig4KnReeoBR1a7JBfkw9RBsZkjBFvUP+7jrAXQ8uc2ScOpPIZYFHAjR7OBx1YFCgd
E3HJKU4q9ymZkaAN659CGo/a6nIpwgvmqyyPR/L0Ra9n5jUauX83clkWYGmYw6wsc6e98i+b+2dQ
nS8jj3iS8kEE4l6xEcmbBEAlrf8HJYVydk4fDMzAgSdvxSMB+YnLJL7QRmTsHV9ZHy/MfhwGd6qq
fvnH5ZYZRE5rTJrDotaUWhnSrJe0m49FyPC8euhFBKZc2RYqQHsy6kaU90JCD4jlS9IbCWt5UquK
FBXqdEypoKVKtncVfqTJRBDY7boZM0UVhfYCAr5GQfQv0l95IoF0C2YRDC4xN/Fa2RBe7nkk9/p5
LiFWSWXfEEipHY1Jk1jFioTRNmghN9Ac+ed/+bb1O/e1F4KSbg/6mTBQ/4nA5QPeKmLHdIEGNUGN
IXBn9OpwQxFiG52YewGg02XxbLepxE0TKlw3jOrP7JUUHIqZUcKg4B3VUM0rVQSmTIeqsCDVda+/
4ZPagLBi9vAvHo4+7pffK3Jw4d7Pk5WVnmhBCPkXP4P2KOHlA9VbQb/MtNxvhmUxJIhZO/yG3KAL
GzoKtBq4d5oGOP8ByHYtftnvEQHl886JbxRT9kiw9iiLVNa/BvXXr/hSOcEJspovbLncKFGgOYeY
/gAT+IqFJgKJPwzIRoIuZXBKTvdb8fh+1UqhMn7TocR3DJWd3+W6O5u6MucqC8hMo6eEEcmyHKeo
yR1nZiB2K03Qg+I3d+SNzMb3V2lMTHFVZtPq9JcV0P6FiL5ePrJjkxNNrp6TQmGt5AbplwO04cic
PdgwIfbe/DgEXEZIx70vPSC/nPVxgUkOG1LU9GxgULhEPXT2oSOlWjdLdY1zXLnLoK+kdjvr0z7H
OLopjrSujes+OGXpclc9zJ2piQ/TrJ3Yh3EWlGgQ1BPMVmgfqijIjRN5Nwc0yZk1JCI72+MCCZaV
6FWTuKm8Im7EW2Cld/buJxsiQ0S46KKLwR4oqHChODC+B/+tZ/JMDdWJm20Pnva150TC/F64A2Ht
lnYeOAG9tZa4gBu9YZD82+K/xGobAPkhaK+jFf3WcWbVp0+/NQnaeKmfbMrvm1iKaQuHvmKhmAU8
m5LL6YT9KzjwmLlq72jc1qsSiygCADHnJ2Fu06JzXlce7/swHLTHEbipE2OzreEIDs16uHqlAv/0
Sb66s7jp1ay/8NjxEqh9z69gcitek5fFFqtFYkGgs+GMgeB1YQBV0okOsf7XBEJ9VH6DtVwV7RAU
yiEe+m7cPXm9ggsS+M5/dLo3lELIHg4MwL1kOHHGz8/1957dX3JCb88QKN2RHu88bNC2di42KrmV
drj92tNt/sFMLE6zxZAdBAGqaJOUXXSdKTVxThtqbKKCft4E4hhjHzsypPFf2aAr51mvrfVjkN/h
jOe7LxiHrpPs/3dpgpInfyi5it94JSuaUDSYi5T4+ZgilTarZdo/kk6geR7D9fcwBU/M8D7/MAuC
wOXmjZ6aT5aq27zugVITLAc4MuX8mhYs1HTj0IVNrOTv7JKMvinZTPHHdJ016dg1cryRAdUfFLXI
nByShfQwJwNVwvoTE2RN/r7sw3iIR8rYea45q37wjb3BUyT1kXJiTt0VwyAXIgeX/fixlg0gsqzR
jbsSJOiwEMA1J7Tb7IjBYMkNGXZIaB1GyLozqjRsH/Ww8qqjlw4FBwArFNZGBf53r7yXKhB7PZTI
QFcAasAEaQI6fU0uqkLV6oVWZ35nonM84V6D6jG98XQev3vgAtHKLyR3Uc2LGfyrniiQTDEEkHNj
Lj+CNslRRLXTdMTQ/jFJIz3lOerDeC3veMqlrFtmwmbOiH3SVQwgo38rIfqgydOROw/Tx+yfvo/U
Dg2QuMK9Up3KuuSzFxXEFnJSUTpHSJu5Jz6+dgd+nN8avj6Q892EjycMBKfS3WsJNjlWVRhQ3ips
8h6EQJOCs3dyCynTj4pMereecODuc6D1nxLu6LozGyYSKMq/A9WUavlcWUepw3RmrTWmXqlGKgoN
c3CA7pmrz019kgBle7Vp/iXndpEkNPIoUZi4EiM59C0OhIT8DtSGktycFwMaw/4TXzrhWx1opv5v
S2TMG4xffgU0BDsoNkP4F+3GMAeYE/wAbmx8oEMOhAaBVdXwfsw5zfoR7JGK5Agj1W1HGfMsZmhY
y2R4lCFSqzgpP/rRIXW0yTxX/61Rv2vSCgruUs+DpaEK8cX0Osp3xq+G25Xi7md97MYIwlL4Hsch
wQKP4nv2KMfOfaGElVMVAbTEOGC/p8a5QXRXHQRQqJ+k0iauQFbZv5KQdjhqRiDcnkGH3302QuGa
AdmoEiKbzk1HcQheZESppppno+YHI0KfqxFu/+3pwcWKIjoEq7S2xP5I6BVa8j6Qra8xrSkDYM4J
AkelMzUWpDKXstmVyio5cHC1vRwFNrPPj+cyt1XTByzNPNxRt4pGzOwDWYJ0BnJOSRMx5uaLPRvU
a4b5UPIK8EEj7AK9TabHnslpdVVhC+l3/LN1mJ1gUSM+RGXRqrPCJ64N5EOwclX7OymaUFbV8wPo
zVqIxYMMYeki5nXHX/UAoTgsQ4mrrn4c1iCpWOYrWYNiYaKCVK2lDZPhgICD729apRfgO/AX7zgd
5iZIRi8/xR5hJqKYzB34rV5qGI9ezLnss9zSngsHmeL4Kdnb0tT5WBVccQLZcTFDvRu7ZuySmLAy
XKvWT2JoYCs2yYapXXK149un9rOCT+LHPvFG2Xt6PB4Kp982+CofEwCvd59iP73bsj24Nrfx2L2s
4/0LYWYtMtRS40exdH7fJdA83r3aRsx7yDy/3K0DRLGc8lh1GUtlOi2igMJ7tf8oU/LntHQni9L3
v23/yfE7cbOl6nC0UaR4PhPqW9aBxywjyxBF9Cls268bpH7taMUg30Or0hmW9mgzhKvekxyKxp8F
oXNerZaKm/gintWgkt/rzf3+h69nar9gzy/jMFfx9u9Et/bBbFzf3XqVedB7DYHayML6+doYWeJP
4QVHcB97QASLj3tKwT3asOW1rZI3dXEkmbvygmvn0O5589Mn4KlIWhSiy3ByQ6Nr/xo/BOFL1NcN
8vz2OZvhsGFmTbZKRdJXsn/VikOnK6EA6lsuktvIpJsLmyfBzIBSwvHoZzoah+SKij8RSh/P7MfP
9VCWQ68CEZxmTW9W0nT1nmPDmYyY1P/NPowtCQMlWFE3FM1R5OEMV2Wg4J8le9fI9YR/7lHfI/zv
1cIJM7D4bZLWfgCwfnbIDzJ5fH4O3ky6zF3ERNT81Szqu3/dp/yZ7tfWtg2/7TjG2V5bgT1jVtMg
mrREH70+b0PUdARh6zSjLvys7JHAVDHCClUr8Vla1aYpZfNRiOoiAlMY3xLwOcOCfuGDC2R9t3LD
bM8QQWYmLnxOxEAUEDIuFhYpRWjr9zVs/BX3gqFC2etc9jdpDBwsYs58xlUDHV+MMzya+Ls6crUx
Gc0r5OGnON8P5HyZ32pHn1XysdxPUv8f8v5iCXpmAXhhczgsjGmcONaOs9lOOpLwD3WO/604rY2T
keEyHFxI4AfCFx9b9qkxNpgAMbvEwqApYzQ/nIFOeAZHFYbJMhfXypighI3KhVARnQ39ifUvh3t9
x5QL5VQ6A2/jliMQsbNIbRY3V1KsLNVJsoT3UzwrcMTmRAKpC3fruwV+IyFt7iHDsnYwASxjkTxe
H21qAPUGtGIIbZI8V5of+cBV0cUXS4hrxTw6Ixp3Sm/R/gK4UyMqcHK4xgJALyHEexTMRifg8K3n
GaFdgTYe/dNjm9UmSb3OVjd7hcypaCRcUf4Mqo+JkqAQocNd3zl3JZwxO9YLY2QxmE1JfSUr5TqN
AGRfoPP3K4wl8ncwPAo933rH7uCrAws217R4gegXX/3f+OhlZA6vAu8jQhSuU9gMM9BNH8SAUH+r
Cqaqg2DVtqA2zXbS1H3x3m3eixRZt8LP9A2mKUIcnPTlOQJDF4CuENFF+fqCEMJBC9OxQtsGAlLg
vk3djVRIECXXR2wGTVc5UpoWbMET7oYJNzv0pXx7m+ZoStDZUFKn8rglsGavpfrqV4cg8zyDBmtT
N40+5KXsf+2DzoC0TlcAHE9oSr4pUgL1Ms46YNHItA/M6BAhF3svTM12QOraPn72jSlNNGzPuXkr
uRYO7mo8lHosT652+FDKFuCc3VYkJMAVGdwwFj/B00zu8wOm8fxXaw14aFeLdqtodjt6ZJh6hKWO
Fi/nVbX0poltDPjwbIKiuFR8ggo8He7dLcPwWWdn1VqSiKtrXAwIozS7XThUHLOv5onLbufsZ/EI
j+jTz1ANUjSdDNWxZ/44ECgIR51eKhdwtXVIG68dfnbq1jZLl06ZmYoV5b0y8V6vIyn3g2vHoHKY
rktf3bbdpy6omOTJuPbf/38Wsx+ICipynMYnHi80rw8gfoYPuAmZgG/wUsKPzlz3WRpPvKzIm58N
OTGhrbmL2KqJu0gD+a33iE7Ah8LJos+S4sLkshV3LmU7UshhOiqnXscs5HYjcX/9hxQq6NVHKCJT
jpoZ7tkPsu55n953r/Om7TnABCw0PIyZwd73eZ/FDbuEyYMC6U6FPqee9aI+zBZ6NTgneVv5V4Zo
/hMT8jT+gycSnKNCXPOm7hTtWve2VCf6DHZtrXEtIMLj7zxLCLNVBIMjZ1aRRi8rCbK5FxHBsEVl
x3UCHMBI3d0v8Tl9xuEw4u+d1kkYhBXwt8uxHhh4BuoFXNprOiMgmEfsie3E2TmcFiG73oJfb1WK
S2XvLU8WPBXfwC4HMegN4kHuj1/z2as/DHgE93iCJ4fVTXUFldkxQ8zp0du3HWw+h789575iG5Cr
/kKjBXDzOeqUx+pM/7jOO2D8iDkdOp5+0rA6dIqyJOL3tVvEwPTk/5+mMuZTAKBKDhC1tHaayEpF
iC8hGsTx/Wge3iO7p+cFKuLqkRDT4tNbX7QaDWaAreqNRcPsfzXs3j6vs2bdr8QMBIPqr86nLvhs
uaUAXh8aowNiwO9C/X1yh2pBSasAzOOzI21rpVKksJAGt0jL6Kj3lw9POnGsLs6lrNBZtVNHF8wA
cjsH2BMBJXV318GkOzK0vVXyh1LePZusXosYqJFJ4A1yXDkYBliyM/bnfjKIJtINIROTAlqLMvyp
EgFocfQMub52Qv4X+b5lTye4TIejxDiHRds/5VprHmRLxKrPF2REpwvh2YabOl1V9XX8PUZxVgWO
DXhj7Ns3ArdsnXZb+vTidc00UaZmDo0ljhF066bkwIcf7Y7CY/CmsqYnowL8nuon3M7TQRVKXAB0
i8HcOZauDrx+T9leBUd4QzSK99Fh/maXcMV/OjUNNfY1/PUuU/NyH+HYpw0NoIlAF4bLCSWEILG4
VA0EQC+6uxE8s94s8yxII8GgUewvLbMO72OpSddnJtAYC+Oh6mo3WeGYrgm7ljSZUQqBGmt8E7nd
KPdye+ryfZdrgaxQCUi+ZiMZoAL5AT+JuF/0YyazTKJbS7j16pICiENdG0McHBGaSQdVmPyvAukv
WKVZ8A4ZQKehUvqJAvWPr42/hbFQng3mtpedgy+3W9BjTH5ApcLdXnqGFFWzUKNoq36i7Tv8yhf9
B/bvzP+Dj7OQeaV9PHyu1w898+c/4wdKKk53Ds86nlh8nxJS1t42AEvJegqQ5uSTZmKLi8JVncUZ
USoPf4PgSeU4t+GhV48kEU0py1wS6M1D9IzhhNfoONuL2Tlb+7+sOrJFw7CbxJN2m6sB6DwGqm3K
0aM4TI35OQH56ab1hTvWKFv9Onqq5IkyEVp8dNN00wC4qXmR9ufaEqV07uz0lephEY+/h97tWXMe
L1i4lEav+Pq2HEew2C3Aw/QPNOarNIWUZPRI4S8W6HtggFR2oAafcSM7gSlYa2oayBs2zLXFlrBM
cSr+t7HAjGviwtdXAOSjMrxTz9iYd2BaLt4NbSNlnl+4oEYawVD8wNwjXrirepz6byhMBBijfN7Y
Vj8csOJVc2XQ7TW9opYXV9X1x4Pgt5Di6etMfU/VKQQuW5qmhCgtdAo2hTtugpGneJji38I9Z318
yE2+OfXZ0PvudJlOi/SLv8pHHhf5GWWUsuKk0soPgAJmcBbO9dl8GPLl76c7RtRw6oxN+E+eMaJ4
4vX0tweUA9efsqkCq14Bx19nJ92EiMT+4WobKbZc5qmtofiSUYeEcEJu2321Yn2wHRI4X6uGbuZJ
er1SP8HvMz85Gs2LE7Fdlm+4GREyzOiEeGams/OY9t0UvxTxb7rgU9J7kIy3UdMGH0NUwVXqtRIC
TobCFxAH/EbbFd80OFoBESXcx6lGBObacZLMRZKhdoc1Pm4/TjrTssRw41VnkOFhS8co1TWOlevJ
XlVAs2eUZ4li9t45FSX/ai5HuFJqU9oYSNFNT0m2Hs05nvgz62s8opvK6l5r9rN4BEN1eQgIaXCZ
o1CqUpo2shMsmKVYqGnVNxHCzFI4A5TJYuUw2IjbznMmxGhZoiaOtelo8dbGgSJR7og9emXSYMjQ
BHJsuZKs9OJsbTTEY5mHDWZCDOOmTtwIeRaLdVPK/Z268ZZJuZn3QqKBOfT02lgxMQaXsGooIYGX
mLOe7X8QJNq4YIOb/S1NglbouiTnq8cWdrKEqM2U1d2SeNz5ci2OAGNb+OpXv2QyTsdTmCfPF9Hr
ug8kYPCi6frbMUuV8Cx0V9cEAXkTj8+oEf8w59fzSZJ/MnF8TwVDDk0bdUR1vL7wg8DOBVpIG6qp
/JHNfxRLcpO4rLFQeQJ+J1jAgdYAuWYi33CyKSSQFWpNAfGaYbkvHCc85Rd+Pjq0b3UET5lqV6+h
IWqSmWrs47/nroV2ZoFSKRy0KMRbcOJQZizTL4fGAEvEMiAnkUaRUoEX3BYFx94gacpxYlfwbXQH
9kD1wTiXeq0x499vWFhIPCdRi2oWFMCndNgfKONwH+zxiJJZsrEM5dtLDBuPtgRLwI4FRQ+S6T9S
A9eK245UKotaT36ZTOTavwLrZe6G6Eh6SjKGFdEKsDYFcxVdVPVFkrAZ/1HlIscDV5rmZ5xB+BeE
luKPL22T/iNk2Aw9QMlrG11p1L7GhC4TNQMmEBgnIprHVi7vy91GBAu5hYznteCTItZD/HfuwfnI
Z+nGTi/rhN8D6adWRRtP2VaOh9wmkInO+/YjLVLcBddmf42KMiwMTjqxjz8SB/ccmTjBclTzcIfp
+uyvanJi5xyjH3c8+SAxT5aaH2X7Af1eNXTg0y4JmohjmrrPiFMx0HQNF71uODcVch4+aLAPbIrI
czkyg9nRIrcq1I9W4M0zOwvWWQmkBsbNm+c2uFMI4m+qPCAWlwSku0EgT3NO2QaFJ5YEGpI3k0HS
SbM8SCwmFFAg/sCcsT++vxcsOrKzHQlX2bW+lWatvMyUOoFarcc0jxT4q8EjTDLCdk2eRcrOfMW9
FryjcjA9pNgZUHTEMsWyB26C6CNcaBOMVLoY7weUkyJRq9yxWConQlfnQhTQE5IOaZT6BRg7aZtx
RLiD6gMU9nhiwksjYTNcdJ7qx725m34hTZSRVDng3+1TdfX6Y2rOz3M58ZKapA8L6igode7t1jLe
xmACEsNJjxrEywf2fkOeZU5YDFs/9SF3LlyboJOfLLfD1x1jvNKm6f2+OECIEOm3fTdWKRsZrzZP
CvP0iwX55aI6eIYfuO+3buDvPhqnLWjLOHlxXbv7dF7vW7Uwezf3JAKbuBVpZ8QGe8W6PV6PEuVC
F23fESPHesTa7SU1AuPDZxDnsiV97U16ihoYpdF5FtVOEgaQ7G5iMBjNsUPWZ6CjsgEiQpa6HGhX
Fwj00AI3lzS/gZFkLaCRi/MUpoPi1CM2NY794RU8F4X5qSyy3CKfXnfg+cWm/kjEG8GPl56DcZL1
vxqElFyRk5WfbbN+8aOR48Wb/yH/OSpVBW8ThzNg2nuWrNdhk2Wgb035uObohrDej50liG0YbP7a
Lbl9jA5GmkOiW/NYyBn78uTH3Vfbw5AkN/Q8vUClraym6Hs+c/05Vidp482bvVugwXUZrf80WzZ9
ftSmjAJBfpu1DvzHv0fZhIejtYjA97LCvEKJgIVQKq7S44iGPnDiwgI9KbYrDpODG2sGfMJ6PZoq
kZJjmgM3zzfA5d/56MXGVOjFnpbreSPkiqZelvKGP8nOr0z1MIIqlwkN3MyniXp2gvRHGDuN6ZHv
0HdJnIwg2hxlxYaBLCfrGn4n2ENfOX/qWjYjMzuzsuUlZ/2ETCM9Man/kEsAa3FoFpLl0CX3NHQs
CqBoSoLsy5pjUuswBtRN2UZZjX9AYhbwNW6jUrLuYBzvcbAqsaDutNvVfOn3pqQ5JQbaCCxT7phb
CBFgPLUyrCuru4qd6PPXT4LD9oCJJxFjI772Ha20C7QcbzvGMp0+kW8ZA3pWa2EIxUIeccqpTBYC
VwlGe49CjDrRxe34oiar08Wx0zW7zygUsJKaQvSC5TDiNGNXScSufnF96P4+bki7wEuPsv84bfwm
+fyUTyeUq94ZB5On8uhOHUjrAKg8aJdXIGfJFgYDzinObn8qYv71LjS+wu78Gqpl24HGVo70f9tl
CUOnTXIEIZp8j8WFswxDgqWJLMIxKJgduIegL0voRQ5tZVYBepwa9ZjbM4gi/a5k0R9RaYuUvEya
RHK4x7g9WWiyUEewQj+mMi/tKh9UWsm5RYbCrYqXzzNFqcggyUKzHHLLEuhOWWj/YUptUN51hSuu
f8bCsRTRM2wyMX7VvTYhFGYkf88tbEEGrfIxF6VYZ1muN2B+4nvpSd9FA+FdeLUC9Bj3tZeCjMke
5CrXPjYA1NaFu3ZYF9DKoIiojIsbHlfwCQml2mQPYGaaHlx3s+BAS6gkVhPzXRpk/MbcBuQ0ZFdN
Oys1F97yvCFeYleP+5pH0I/E2UKVnVyJq204v1BK3zkTR26qRAuwsKxCrtVRpzuBdnaTsObudXH2
yMhEeccKQQRNt1SevM0Z3CwSxpC1jv7X0Bx6Yqnj+L04cUYCSjvoU0TYWS9RK8DW3vRCd13Hr+3C
3XExJFPwf9jrSirWasctjlH9RHs/fZFSYwbKwhGAG3WYnXyc/x3D1IE9ajVOh683Lat5wiygRBX2
lKWzkiGXFMIH/ehYag38qcQAFZ5Rfh/eV91CdBQIccZdB31Pb81jY69z4G4KTsF8+ZgOi1Spq2+N
UAED3H8He5djipH8yJP5AbpxZKHWCoZp7ap3NtCKoDYyb7O/hRR4sIH15RmsF7SniWQHyR/a7hU6
ybHEyNeBZ4ISrogZ9pRSoVDHQpJc4TJ+24GdoD5PjF2ConyphrF9YK8JmQZe/Rlxg2ZWymyEPrPr
Muj5v0uTbRSHa0BCUYJQ9rw8TfENc8aHhgHyyC1jTdo+AXWdYU8YuN5RJiO6XcSgBguFwAxw6H6z
L3Aa8nGrgDvaHb9t2bIIb+MZtVovri/0CnW2iAZtbrTQPJSDuhmG5t0++NRysBUbNKsgAGM03vhC
0MZEa+eX3L/40jX8ygnYrhTChThq+PLncF37YrCdQQCbZ8I3wS6Kv7Ah9qzPzSq+2f4nMVD5Vwh9
S3yCpkTIfSWOHa5c6eOBZ2BDdFjqWkUKj0RaafZ9Vw7cEdDZxs8siKfNPmuN9IWhXKdEcyBzfQA1
Ki2WLEucnEYmUuQ+jtmh4QgaBtko/5EuMIX82fkr5Cxp3FEQ3E4Yh/se9FD+zHA9+EX+wlYgjtEZ
Guc1CDtf3hFDQDKnclwe+8sB93YrMWfefijl7Qix7fIQ/ROwzXP8aXBORCMUqylCdFAn+9mW5Qfu
PYbxvZsnIY2gy0CZxGqMQhy0Q885lC5PmdCTyxs9Oz9fet8YpvW0IEY/QTAcKJCYLB1KQUcMEJfD
GCF04wiyVHNuYsYC8uXDxm34+d4LjFWcKaUO2WTnSIO9/Eya9Rkgxsi9MzmEvlOu89+VZ6suVyHS
VbXSDmHMFWqhKHOeIiDN8PbeYW5mQQOrYn7brgyxmPKf2uWljv6ksQJ2IrYTQoXu2vougemVqxP9
blVNujx9g9R8AZaQQ4/6ZeveZLL4+ND9CwKYcKoWYjI1oBPbVP8yXYvz5w/K7PssiCi6dHAmS8y9
i3ldHocAQvNe/7Ci4o0BRSk/QFrG92n0P3YKaowyGRJBNJaHFjZ/KdMZ5k0LuAmE3K5PX0W26Dlj
Pxt2bdCs/77CFqJ6O1jFm0OwIuHyqfjnvrwzL7SsPzG0vD8+tZQcsxauhPVxtB8McsrJik52DgJT
iLi9kKaUReek0pZrl+87KwGMc9CLS/vj3UMbe3BtgjSVoCOcJLYc5rArqCrF05FEwWYk4SvlZ6BD
5XN2Fj1qcpUE5OopiQTdWzxkRJmX6peyD4nv1mWdkOkmFxt+fd1vJQ4li6txYlHgr5KXzP3TF5YU
bs7m7Yh8/v3IhI3NIJO3ZwBoO14GOCuZNN7qLqzDM6ojTHwWrnlorLuqTTcNxtqZuunkLwKt+Pc4
/7xUhhrYqc9sTSABY1jy6ia8QYfFeEPMm5NsJZ5cJZWlUYnYiVuOvkfYt28g/6JGHRatOf5Ck1xb
avlLOra5iE0vVEcOH/MXbbNmwEe64UszIc/LE+Hz8NwvBIMnRqimnEq0mcTSWafkQY1MNrZnr7m+
3ezNNbCIdQr9iM214T9zqzXGc6xt8Tg5PuRcJs/HXGAMUgWvZIloyqsblj6EHCMc80lPtxZkr/BD
u9vvekCCivUmcSZfb3d50U7fM50ow3wdANgpuw7J/j5TL806Qs5QbEI3gAB6MrRYQHi8kVMUeJuL
Frhwmr1grBd3j13I/euayKy3KYpgTPHaO1aLKAzKMFzKUIofW/KHjr26YT8UDUj+slmZamPC7RhR
doDQGKjhbSJ4Wh3wrqPL6cuuyh/7nmXJ1iz6G0LCjl5TpjhPvoic9X/927lJLf3rlhEYWdTQRIhS
/RvffvEvgHAPPIk439J24PUAhwEYjTBghd4e/mG+FnmhMIM33wmS3eZqp+jziWZBfFkZk5auEa/C
Q3VL+suelGwq+shP/z/yIupiPFjffs+A5b8wY2+e5oVRqok/QEviGBUMOgHX/OJX40VFLRGQBP9u
5FNL2oKAsgUGlmYPniba+5D+qFtMmv2Obi0YI5VzNDRjARO9gJtSjQlV+vqMce1nF0EsJJFyg65H
7lii2wgRWZDT7Sdn8r1W/C1Cep9Mspc92yNfKuXqISoS8orJRH/2bvAJV0yD6lBP8/01PXLhi65G
QbM+sCGDGQWXIo1bG9LtzQpvAN1GA/+emH1sGCU+r7pzYzn668dqeIf/+0LNaNfyo5K4tHwetbaR
JAaozfDrSMTsSpdkvhUWFQUattAoiTi69zd+Zg1kNcDTefLvyYtv7P1oblWcIyo009Uq+qVZtiHH
khWaFTUJsB3PSUHRfXTCXThv+vpizbMV2igYmI9A1Iz6LOBaGlIeDl8NpdO0ZbDq4Dd4/5mBIY9B
qTTE82ylXQ8b4MMYSVTHR7U9EA/k1nMfQyQ/6L7GknHZu6QvlEVmFlY4ZzC40KAqyq5coK1PXa+z
nGMSRDUUUr1jG6pyGrxJNdST9k0yO26O7JiQyv6es5SAMSjDcxV26Cfwoa9tAnpVb/jFuP4133Hu
GoHy1NnuLvXAF0ivJqy8hVQm/jcehDzkf3As/6fp7H58ptwIwuTwLNxCY7MKzroqRZ7YlmelHQYD
BTwf2+m6J97H79dBx2b/CeJ5pkhsmvPBpq3xMxf0aTDVK03mq6u0UML2FLxIAs9rvmYiQTUkULiu
aB6n6/7b95ynJCy2kX9shneaL8BA2l1KQKoSNJiIhFB5qZ37JOcGC3tfZapl0nTpafU0ebz1oTVn
TV1h97tZhcH4ISWx2Z312OQdEg2O9RBgnjjbBojVhnLJyo3mwEbHtwovuqRDsWzG1ZUVHuNlWi0W
XsOB1FrBr/+o9y72/DH6ZewPB9RCD8odsLVI1r48+cXoqbj5FZxcT5v8vbzSRC13D096dUs876f3
sCrTmtG5wxD5EBO0yrTzMHrhDZnxGqduZC1f/sOhCdwJ9TY6tssFiFx1lZaJKBvEKJMBH3ZQydTS
Ki5mx3pHYO9AxdThw1Rs42LxCqXL10GAPizVScq4ZBvnx4ERlM3PxrgN1906379rf2s97IJIigPX
zrBmVhQv8WyjkKu7hrT9VD9WmlK1Rb15JpEGtMSUKgdDUfKuAQWKmsxKLpzB3vcZ9RbZGyiTCEXP
eWIfa9sLgnqO5LVzYeaALWPnK+z+sRbUSYRsG5s6kzssYxhyBsu2JdqRv9g99j4+Us0Vbfc+Ge1h
iH3OLBgKjTyO1pe/KJ4yn3jI6IjAAx1l6o2i+0XqVowky91NrjUHkajiZMoZdK6QiTP4bGKl+1XE
USwY/04sP4MMJ34LJEyTtY/KpFBVgWrrMuSijQFpOgsylZ16AVRiFba7qRm9ytRLgqbSsolOZ2SC
+txTyzbIc/GU1GeBJrchA+NNxYV/IpNu5QjHN7GNyxFaaoaPHv1azF6jJVlR9W8iiLztyCGsj3Xx
RzUHywYwKQ1dbh+KSYRYvV5xdZSSsvHOhuCmnvzwDyrN8RHt8Oh5y1ZIdwsRXDpabjMbMWiYNvSp
8DYy4qLHZHHdVUYn4yK8gTJXbSfPxsiKaeJFL7/DgPMBRxV3XoFjlXpdKZjBjptL0wSpjyz+IJ3x
3urEICr2+3KMJi9rwHQLPyww1Pc1OCs/uYYzMtnbdvzfoAYFj1dLms4F8HhC6ujqfXqdhzRYpHW6
3OGNcM74IsgA69ZR8yf4jrfu12pOWbA1Gl8DEPFzZsJPpv2zApsjRGzVnRO+EtkZgww+OngS3Idx
IBM2cu2DBE4+aoQ0WN5yUyNF+GeqjNZCqb2eePgzkxubM1qVSPrxFCF0Gb1DXkV26HLpQTl/LVyR
/P8s5wMx8R919hOVgQ/HX1Jwp6hGXo1tjPzKcnWHGisnSrFGudZW16x5MMlfZ7vfpsxv6bxRMU7e
mb+bcnJH13UL31dOXvLIebQ771tBRzO5zhEpnCMzFHUl6lW5TssNb8ptVxISOd2MbtcRlUxLGOfo
568DNDpbldoVv3ukyHFlN6Z3Ehhx5KabecfsEAFnOCKQuThObyiobYgAoktQVidkSY1Ml31mOxLV
kul+OyroEop3Emo0KWxkdaMai14UnWXHHGkMHEt8ZCrmXC1gk4LQn1OasMlYJ+QxTrE1SjgGpqIc
EgxF7qBz2VNc9wI5offX8NAHugyavqZPWbEy0RHVzGlPU1xa0Wf25DrUHJB9OmX9yil0XbkyLUAN
uqbfGMl1jmI3QbpiSlQViWmkTR+c5ibl9LzK5PLCcwgs6ZZdgIRLog2Z9tlJJS/y4Te6CltqOr1t
ZCajmqH+4MyA2+ToCdvl4B+OcbHAC0EKCLg8NQsPIANNTSvfsJBeA3ITKDT4c5Qho8H3DwQPi56f
lhNF4AmxPYbMDwvk3fxkuJDOfHWUthFWevtGXWi1YaZZsqo751hWiQdEwQS8wVCssQybZ00YgwjE
lRWKzFra5hAspoMW930UPb8hnz92bvgPYGCOX4NBbbwbyBEjmTr/kL9h2C3h+p/31FkH+KcgK2xK
JmjuE9eVwqsctuGwefJuA+pNYOWdKTC6WvAAYOaiKPthNi+zwVEuxtybTLXN5ojt7nFKVfbgVI1H
5eCDM78iptccPC5zyG4ZgJ6Bh09icanqYi6Sz45x+3xZTimB5UZCe1U9rDVIO8fHqGGSkFpv1h/N
hQQqoxjMew3pAEAMKMj/piq97DECPdhQF1HsNUpqrEej9ocLPSk14W/BzqYMtols/T35x5wcQACB
MKK8Jw3AAMMNH5nAQlXjDx5v1B0igP1oXPIXdTzV2W51BqhYXTWAVGcccl2XuEIIIlIY9aSG4e74
AcX+sq4FvyqwlyYt+J3756W3oUSzMtETwqKbeZAleN0iqwWZuc8t/k+A8nb0CWq+jN9owUkjrhJc
1xTidHE9QMcT+WlkjpMPGt7UEFxd1/hXyLlGC1bfD6ERv/Nemq4DvXaDeESd8gHi6xE2qKKnBh7M
+jgN3oV/cY58rk3OSTvbjbPJJ08IH6anO1lBD/WV/dsOCsRycgj5CC2MeOcfiB5NPI5qmmIOJv5y
T109cTF7veBLoBLGbUNkpYtVRy2uu4J3R5AuVnGnu6XOk4HT3kqpfseJvCQ46NWmHWu4zxBVteOU
a/zQ/raL1a2+0ukTrBVP9JWXhW2rnIBphingL0PRfKoobzGzzCQVLGOCnDnURO4uswKX2Bkhx8eB
LtCkzMynYtefNRFN/hAUTGxei9EfzZZDrBnkVoYPGEY4IdYwsrXMeU7wBcm2NOanjvqPzurD+lr6
BotRr+4z3/0PPpt7jPPnTgxiiq8qHeJCmOukRKkJxs8jdmJEEsMX8XlMheQ79kkE36QntI7AMMro
t3E+EZwXarb7AomH5pQ/dsrhLq617lWkB5geFmVJspmlbG9bhFQv7QWLwiT1m+/ZkfM1Rmk7q0By
IhpNmODpTsYwppwKaqQapItdnaInDmIV7qnr4qSGlZDlrs1lrioCTEwk1WFfJmom01JHZZCUltQc
GPHqf1q8hf+i4ajVvyXcpoK1lIc2BiNzvJzyMbDuQV2MAALftlR0Y2VFvbjjvy0pEK6sbgNQe1rn
JSluhzRRbginGg4nzqhqmh5LPP6+cZ4fT9WwaprsswX7b6j7hrKsbWybW4oGVdMS7DdiCKLe3mSL
ClKU1NGze8kdBvds2JBQ2p+vIwIdZ03QxR+iBDac+Oicjei/hbDk8575+kFRY1VHG7Ws/yph4G2P
75ngHNqvuiLeouIuCpRqu32xsu3YbtO2dozimotwFjLclJC/k8ripEi5/gHGg9FwwX9WoMUuqhw4
U4gUzx4Au/2bTCS6UKikUygJRDM=
`protect end_protected
