`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Ugc6FdWL7POZ70z2gd/vtc5vUTk7nmnOc6x6GMUCdUwoDFdT8WnSzjKh5I0Y0m1vniIz2Yp2cAqh
OaEqpXGrhg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FXqM4O8QPotfIimM02hA4j5hZMdmS37+swJBqH+5CsUC4DNKFqjNL9rIKRWsqluRTZsRa8MDaMQ9
jPvlt46L73TR6jBrlzkW28QBwiXeSsIHfXdvFVRQLMopGVaARQ1EGd9/c3iyjwiByAhW1Jt8FinD
dh5clra/xBz77UXR7tE=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g34KQoxuMCd6/UoXGNq1LUw6fACbLJJnWrv+t58R3f0TLzJqS0A/IOV3Ebjdnvg47tFGL0h6wEgk
KkJ8kgWctgN3gtX3NaEq0Toar+sxaw/4PPZrhJbqNrlYzpbn41rhMGt4N8P8flFmXPBnlNDzxaiK
CXCLCtRLBsAS6lTX+M7p5jRs/PxImqwJpXL3sWTQ9/FgY5wwqlMcCzAvD75kTe3CBE3nFu/SSpaZ
jzfpkW/4SpbNqu8flTVbEcex8K/HDAhBdWlBU4tdC1lT4rocPLBCSn24Lr3+Zp16EQgWHu3vbK1O
m6RZFhalcb7cRImMxHmCni7Sit3hqjaHYGNssQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nO6jnd8pbwJfbbg2+95ZO3AVri39Vy7rD5lRj+3/lF84CltWRbtzoUtbhj3ZgpBdioYvcTxGv/i2
8YtJgJDwQkGZm+ewN8eDJrDJvY+jZ3PKD/htPOdIHeirYWvRwzGTlgF9WUelbmOk76/wSMi/zAto
bqrhQOz8dzZ7WRcvgTeX7CXsbfpe6ADgQnVEVq+tb9hzIRP4B0RPAKwN2Tex3z0Mep3oNKQ0SoH8
tBG/IyDtGGYDOgGnnp0kR5vQAW7w4W2OZjMhWVsz2apb1N1PxUQQjRGrB0x4h6RZ2L5Ve9lhM+3U
RqXJ6/P/7ZuTQXiH1fGJhNMUdenwcOfDrZasDA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tUFKsnj0fNStBFWGXviiqLpQAWEhJPNc+y2N668WT4AjUiD6Cfi3MsIoPl3iITeV1NQi+iTF90tk
vvE8RodWQhtaS/b8F+twGWhoCwkNr+s4e9c/uUJjjbM9Gr24C4ej4KKhxPhFNYBy6/eZ3LGaznr6
HLUk5fx8JOSShEoonUHK/qvSZouWlhqK6AzvdFo2fkRAzJHMgFAorMWrkBD55mXFs4t912alyDl/
DfNi0s5x2c+pKbcHCYZNbNjIi4aZsTaqxURHXQRM4slSn1719zZ1oZKGWLz8FM7ZNj+5bqSLWZ3T
iEqvWCzWzhrwP10FIfcytMXWL6XN62+quaWveg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GD7wPrCfjGn4OXkOOgEMsooysuGTy7fuf/t6s6ed8hI6eVO1wiRiTUr8T6TOFMUPz25Fe3+AjAsj
7GJP9S+ylHE9/t8ljSrYjm+tr2qp0pItUQHlfnzD1HDFjcU2GQx71hUggRP7HSTXoX0ZBtdMxJsx
y5wU7l8PME4Z6+rFfWg=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GQnnfXcKvfJGHibasZeBo9w+cQuQQMi0GLH3uU5kRl81aYoMeX41ttSWKNlAw2smlufudIVWIqr4
1XDM2abRB//KO5mDmKgYJIg/tf9731+Bdr1rCZs9mQF4PIroKcKqQa74O8/Yf0vQN0bHupu7hLbR
dvYSfOCD+cuomPjkVm7OlHAeJENPiNxOo8qROXxOi11ob8PnO+tzX4HuTSNWvZM4owOCdeV+bfJu
P4INquk12odtGIE2qfP62zVbUOWXx/QWHOiIBcwofde7bjvBW8FaJHBlvGXfqWCbzuAJnK5HQnoa
ghV+DzALxr2evIF+0yjPKB26Due69DJlFy4fEg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 102192)
`protect data_block
zZ7suY20nTZD+bPQR80LjG+FGwO9dWl+VImLf/x/0fQuKitXs6xGaRNYVT+X3oTpIHxDQzUvJyMl
NNz8Po3IyjN2rn9GE8ZA6MtK657Rn8bm8LFmi50qlZEG5cJXx4BUd1hMyIAoWbG92O7091Tvtnxk
kqSBYewLTWPBLqLy6jjmAn6pIlT86GFxXN0qjnOCjKinDwxyLLaNqR5X9phP0OlY29eY6gUkzWjl
JOoz+PpFNHnBOqrdqVj4jWU9RHsv+Tlmm5Ld7bp0bEnyCA9uIbaa/TR9woCSHMuCt67Y/d9OZRj9
hyiBO85V1QZY4yNv0vfc6OZiL2uOQg1OgqekYksVUZyM3kSNZ4Pm82qPS8cxBLsiDPoLFlK5dp5O
qOv1nqWbHUAaujrDSAS9R6nz5XSCqIXXu/9tARQIWfcoJYudwEFyS8sj5HB1LIHNfF+S1CF5Q8wH
qTkWMevBOipirtZlxCQxh9EGm4FUECCGabEF2ygWSws0xMZ1lZ17P3WplWZzvbMcmni4DO4E214u
E3PMI13SoFocYl96NfGIS4oVQ2tLivOMutm5hUql4pqvtD+Lqy18/ceh2UVEtYIo8+Ey12+5bFIh
s83xESERktsaIlDI2ursYugJ8Wk91GWbGM6GB/UJnq6mVjUU4ZsYvDnVZ9ylE0NtKwOUjz3gZZk6
iYOL47gsvppR7QEGdJSQUUiZhVfHpaML9O+fb5hECbEUtM/jIWAr4fk2bAOadkRS/MPArN23iNc2
+p0ge7YQKBOLwSZFQZ+7A5/uw2glGER9CDx2jZZIi0jatw+YM8btcLm9uzCpKvl26r5rfMtf3ggq
CQyo7PsmWQkrLrpDqh0lUcnf7MW0+2WqIMVrMyGHoo8QEyzyIouIao7XI/AG0qudvE53rzQe7Vtg
0Hnj+/R/a7fhrPhrOTOgbS0yMdJftUxWTKqOgQDJyyXAFhZhHhZZL8w6D0lEVe/YtVRaBMOm6Gl2
vLA9AyF4yk1gRNw7km3aD483GfR8gUxadaFWUussBRbk+jnnktaAUzyUXZdF3QT2RGDdd9ZFVy+D
iapYgyv7MxOwR2SAlRV4du11tMhu2SPmUsNmnmvEmWhHsQXRoR5SDEwLPnLOCWpAWj9Yx4Vnp6C1
DuIn42MNb3uwEjy/RbxCrmWVk7BbJ8yg7PYw1PUCEWi0YJzzODxmOwgg3XcGYdJ5waxfFdECSZIi
AZ5EMQ7Q5vWLgo1L0TRWXi6FOjAks5xkh2PSV8oU0NjFuVnksZW7ZZGrREE+EN8YXRDJPoU0n/jY
uKE0tmuy1+F2fEzts0FNq/Wgh4bwkFnVxvFHU1CQGh8n+MD/Xo3UEKpIg/PQ7FJ4QpmkPtdcsuST
Td0WsvDGYbFdWX095VGcG6ApUlrKZHXMfz5mH0DiDbWkz+jiL28E9/rx4nHh425J2ScwA3zZeuup
M6//Qtf2Qub8T9JmPAzK8zYctYap9BOQtK/AzB+UEWC3OAF3kgSDxRqYmWGXpZXnEhvczTol7fso
F9IVgNJ0s0b/SuWYdzX3owkoOIl/5VnDTFZ4k9Ow1QTY8QYVz+l1hTBeOHD5doRri48ZMV9aGM37
gcH8SQWeEO/nDmBSqdajFhEzcLJNkZpIJzsGh5B+IEO2eDYaljjotVYwFDyMDGdKpGDVHuvr3d3D
v/1tCGVVwiP3G2E9Z4tPjYUy+FWNZr4gh4w4nGXcohdhLoCj1/JvOcxB0khcjSR5OR0PDcJNj8rq
ITy4pu7+GNFE7vcy2MSpHrz08hZ6jTWSXqfe+GAc91o9atTIQgKUxVKu5mU9L50I3g5aI45B4QaM
FS2so+GuoVyEANTvmYEsRKDt2LFsmtA/pHgo906o8REqX/SiaY5+Z9GpBwP0gayXZ4csHQmawA0s
Ci/MKtHjVp4rendWcz6I3Uu0H7wOs8gVbY9yZc9KXZgRXrhtb529EaSptb1s8ej7ca1Qrdcpk8Dy
m5Jw1d/n3FzYePnew8YNnHuNnmlCuNLPqLWMtlzUKQ75TazWp2PM0Yl7RSmdPMkHTQ5BXnSLIuQa
rk5JDVyIo3OV+wydl8ZLVhaqjVn8ZRRfQuuw9xtd4r5/TJGUeSl4/5swFjaQTmSC438135+xJmsR
cA42DwmlmT68eKNjBbyv/LLVWHV64CBCKnHAHe7B44Db2XYtAduZR4saVw7UPyESe1t3rOtS1Sg9
6FP91K5JMEfUyCF4rp9R//VsJiH1e91LmHqdCsczVZmIyB5Xd6/WwsYZc0ZSLpupDqHmvX4MDFjr
hnvQmq2jpMqSA7LSUvJ4O3Nhxyc05719su4QuSKA1TArSxeuBgRK2aHauHQhiM5EYCmqrYXtBn5e
+WoCGl7JUEugG37gkJ+S/FqCPHys+wJxDdWGXXULo8QMSdRqN8d131EkwITn0Ojyg56HhdwVSw+M
jq3Ch9nRUcM6kaftU1UOMkimdWuB6MviSqonhHlTiYBvCErR8fGQXuTKGaKEoRc6hjjU5+9k8Cl/
iLNdg0Xrm0iNEF7coqMiBHEB8UbqHZSK+/ri4QC76lPm7g2fpSlarhKqSTrvPWESEOA5Cy923Cgm
h99wPp2PIluFFZY9tHg2UUwSVKdefpa4LsCV+4IOg2bK+/WRo16f4IzJEqEj9u7eHPBfgpuaxuO5
RzQQcOzNFHss6CT1gKgyGxJcxcFLvnvCEsm1ceom7BD/YwwuZt/zWKlFXXfCzh5NxNC0YyY6OIRt
DTkBypMeBLITYKT2Fwswzoi0EMiVsPFhNBdBmrIFSq6UHfW6kBeyZPnUkJcmpxkrEkPhfIrfNaHH
W0MqPXcJZXgg5RyfYDmLIJodCh0odBCLf8pLnCiU4IVykt9CHFwuoveufH84iWt6Z92kqROeeWeb
f2zuyyiOlxsIi1B1xeSa5q0A1t1fZLtaiAIaLalQ7WcaH+kIPeJ+0iopPZrmlIVu12eLQvfUi0pc
LH0vPYPVWIUOTYXVfZzimStdQ97m4wxCxQMd0xL3+NhpeSPDEtMZk0BxpIwKDuKaA/Hen0JgxgRI
QuMGKPN+4oAVoNczsbfyaap5NT3UPLjkTyVDt6V7RZLHom7KPwkloWYtQkJROgk6wVOMt31qyjUf
ANtsi8B83yMCERh7M87T44VhoaMbtHS2m3AYGMw8Gux6oqv/NFpMchKGKjftxAy6Mgvew0woPsTQ
HZdumPyyKlPLHsgsaudBXZoH1qwEF8Bo5bEpATNjP/HV3PjEVuO6G9T8+KJxh5wUV9C3VtVYjuiS
3CTCD9TIeJo6DcSWkwcT7HsuZpo9Jg4+N7Wkx/WySiLpzm4thxhskR7asGr5C72xoYUdO49Owcn5
PycLaN/Q9ZDifYmROd+A1TNVsgkJvDDKwI+Ok5nc+xcNwpK0dsu//HjJfoRWgh8D4eR4Iu17QucW
Wa+2NuiNbfRxOp4s5ukYhHnpGeNBi6yN9FXFYK1UMIErCyK2+OPRf7L53WQmYuX4U5Z4erl7VMuy
VBIVXGmN79dMkZxUl3JJJukBdBN+3XIQHz+RwMCaEdLEhWnLcTMuJUyEjA3h8BYEyX+suWsAd4MY
kGfHApBvf7t2IQl9NLCJhmRXlbOLSSqGvwQn3uA85t1FhmQ4cSfy2ZUZYYaohO4t5Av+0HyxmWZX
8VRdzh2xwU1JxCEBa2yOSKO1Cp9bF232p/YndXiMHqaJ/ZyGUo3qSQDZdGb3Zr0N8gRR7x3cmStF
znyQURV7r/IKck74y7X1TSwBiSoFBFX46tV7tAtlRlecylIk69n/eQwSATtP0HGCt9WPuBh8RNQw
/Nalh3L6zyni9KeBn5G+gO+/aDh68bRfDoMnhNPXj4unb7fDfxJLEYwciSNDRKaIuESZPi3KIOp0
ngkWSJbCeeFoxumtZJIr+A+rURxjaCWGezeTTIulCWJlnuFUMa0Frgxy9y7rQccM8gSJvl1Q70oP
tmMs3GAqxkZ5cl8wzcG3E5an0ADgVRjOKQyOXn2MGEXVlmxyvzHhs7PYIxNbvA3d/wKWGIqPUMRZ
ImXDy5t61TAeYdalxynvpqChB5iKjtgNYIbd++TrqGBBpprU+qPB+hd7nOF4iDMlx8V51qtMhSwF
l87Gpa2FOfQNOfxwQJES6mxTaQe2kxXQW7bfZNX15gUZ09pnLfQZGWsarAV43oa+Be/XQAIQQVlt
SsyRno6DzTKc4vSSNobTF2CFDANhqbk0Dm9Jv8twAtylxeH+Td89T9IQ7UbIz34T9xwLmKsnOnxL
3zAFZwqRSdPrfRFu/SF1y2soWuF3hU1qvONApu5XMoQCCuOWQjtpnvEFsGgmlyxoGPbLOiqUcatA
DQjGKQxHZiGf1M6JcjHc0Gl2L8AvXS+NGZRbtdDWOy7rrakrqcJ1h8HqtZJAigKCy6Ixgky85xJo
rT5GaD2wRqcPgzxnHl9Je4LES1b9ufF8aiHMV7YlFYjoBLxeYq/SaLtKWGrEh7vY+BZqzTaauGju
oEcSOoLTmUKTgTdPcgfyEzzvme+1uMDTQeW893ufqfmSMael5Em+oQ11OBsQjn+xI+/ZNQUDrjTz
GhTCzLJn2x6/i37AO8aA/dmkzzKwykmheUeLfJMCl1UrbaSxRJNHGXw7OPsXYWi95c+QSe7eUWeH
qTuT+o4XbcQdx3X18EsZejt5y28PvotmSAM8Lyg1na1RJH7df1ipiY8asi/eNG0e42YwcXducnyy
neK9JaFLNMU20Y1YRHC1wKxu6Nzr0poGSwwu0FA/D32YGvHiwOjtCNwD4yDVAiYXAmoKZnfwLKRS
4nidCT1yCg7wUhWI1u5+bfVej9rf/o1sM9e2EUdoY3/MBOELN25Jx7dxOTMvPSuzN6GtZv4RFPyA
obHrR35lnIXS3xpoTzZYP6MQA5bZ38WeV3zbwBizq3vl7JO9xN+As24vEtn4FOz/xjFx2RS/0Ss7
ZTAwCCKIIDYNNoTngDmm2/YYWvzC20LL2Gh7QRtIORH8gpICxjV4uRLtZk7qeXWxqi2K4yxgid/F
qDTcLfNzcvxyfrJv+jaM7QOFHPysOiR1xRza1cZYGDUs/V4/KbYX4TVBhRUFrc1lZR8cniJ/aAbV
03tYG0GPOt6p0hJGHJqjmkGYAzjQS72hikoOY5NU8UMMJTrBanVTAz2EIzhUFysVfTOfEkTZ8d54
afjIZDmQj+czLywmixB7krMguZH2a11X9TD+ZT43rhw2zxh9ezV+fx+E20W1JZQQ82Up+f3rbcY5
gqB3gJPQt8kpzPmdQtDyFHEd1e0HhHXuQCr/SSYoudy/jDUZMQ4b+pBuUhtoDA/sNP+Ru5zGBZf1
aqja69LzIojO2NtMSyZ2FMxz/DYnhE0DfZubS3Pp8HL2POucDz8Oj74j3h5uLWX0+cgO5H++o5ed
YlNbsXoAuJkZUlPJMtbaKDSXEwkQ2lZaH+sjDm3Lo+m2TBl/Du1GGMZd1SPK30ejxkB7U1kqPcHu
APTZFWd3dOleyYDW7kINHHZXPiAamDh0K9V0tUvErv9+NxoYOEl7hZMhmKtWtvnqg/2jWPnoihbl
xDixsQG8FbBRNsTx4u+BYtQgGKigj4uDDAc/+FFHXbqpqMdsjGPlwW6om5d/fvpA0djbkIg6i3ww
4InwHaiqhAjSta1ZPICAxdgr5xM6Npb4VAhmaouQyR49aBtEZFzkah5Qb9MRUnLtsTR0RMTZNvd8
A1KxIdUjYswI68MfVz5IVc5WnHHb5Vt+tPKxyRwC1dobGiwZM/X/czErJ1JscSKw8bXOZCAY7WHB
eFbt4dgD609szSBAiDrNTDYCB9eEbwwK8DJyNazELoCyzGpd7mS3FGaosLBkTWSjlSXE6Zyj118M
KnDmqAydFa3Z/SWWGYpuTksGAWDEonAMT68V8OWWrIUzymXJg2BkTMJhKMvRrOKpAMbwrRSWlgko
JsGKNtlF0fTOwH6Iq1+5BG0pQDD1B7KZv4TxbDEUIDC8k5fii8iTpc++gEUs0zXcnh75zfpxXWkz
Uj2N97TEFhtVvg98Oi6N/LxaTJu3out1/Gc1aBAD6Xe1CExXqCxE9eKWVl1c90e2d8tK/Ssd4c/0
9NttUnuBpUWXnHlJBHzXB8E+w7DV6hd5S4gXi6R8jhyeE2XXJUVHHNnIMRQI7J4pXWGhJg1mu2r3
7Gcp+oD9AMHtjRvxgNTKXJicD3qqccGwhbQGYYpcLphM4c1eGrS0FK8WHNKKmDQxUAwFN1zEJLh+
/omk2eUEGfaEJB0rYfiHvqNtJ+4blKK0f4q0rLw3/Tujb+QFGU5dEJZmugvDmjxwN3GtGZc6CheW
Wdlz7MIHXyETm3MrgQvUC2J8TLGtKUzH+5umr70J6phWcVypOmw0KdmZPpl4I3xqUlh4OMueKJUs
L80+23Zsnzzj3CyQRTXuXKLmmbu20MGE5qLJTZE3jxKNh+lArnBl1WkDzHB6/+YVLxSJj6kTSbzg
Y3bl4Lksx7sTP39Zn9OYiTE0T6R7Vh1ZU4yne/nw9IhN4NZtmigE6pB8EtvjANKPTd5m3uju+DqO
att2pdCSvn6tw02/3rasWBS4Ze4NLpGYMuIH1J/eAUCBEr7OTrlrZMKDmyl2aKwLrUsv6kK0VfYe
t7OFyQ4aJpL5RefpBClpQJRzrHRhjBLHmShKzLn71MaWdYaDOMzzJnSBBUxu/CrsR8QEYElq1LDt
qZ3NbqM+KYXPD/o0RrElacKFKdcnV3pev4srpbRZcdXW6maZNrqu83hl1titl71TPJPktX/HeDHr
39kn+J3k14ke1CV4mHmrhcRPYNRDKkuzhSg/hdW6ZXBijr5snCnLpL5YMVuyKqnnT0LAnZ0BNySf
s6kxlvjHIaUQTmUjpPwIoVXtT0uoVnE6WB4dhwuDb+oyVRE4xOhlFEyL+Q0lDz42GZTvxk1Sh/rt
t2LeJxnZglhSEsawc4SxVLHSCemPO1RTrQRUahUmvUJ9S0GbwQlDZ09qqz79+8O7VBP8hCemJR5b
mpZJH22Jf8XFTEV7v4UoAGlb8bJwW65m/6Ny9mU/fPpNxoh2l+mu/xOr8bv2NyOASoa33a5gYMmc
PsAo5uBJYtc2yRYniR3zazqQOyuZW+GhQ4F/POYbBl7pXGPoY40cVKVXFGk9HNWnlFJ0xkWKJKNG
VO1olbLAmFEf0Vj4lQH8Z/yR3stLOtmGYD4n5STlZmOngdtYK25cm5uolLkWZfm3Ba2/OvwLEyYv
xyw7LNL6ZNZPUrrzTrZDNeCAKtcVOAmaDQr2WYKZN2I6eEC85K4AavIbGcaQPHdK+x1dqxDuRRQ9
OcNdDT20KT43m3hbofty3tbHiZW6UHOtAF4P12t7GgI1+GRL2Ky7n4kGjcMBrWMNI4Du7w0vY6LF
fBHeS8TfP/joavx163qF3lN33j66IRorN1olMH/FGGYBCFx8DRHK4L3xckh3ncc8KTb8vUR8vcoE
5664Ln3mJSNTzxAxByZyhb7dCBNhgrG8cjuBppvUZ0P/JG9NM308bk15DWSMCBYi8V9lRShRXh9u
qhHLbYpuVSSBi3ZMpPe4XOyVTJdGgqae+rWmZIS5wJCWnZwLUio8miHp7NtXyybhwsK7OKkpnbVh
HdCEtMEkaD2F/YDaG+tPwSiEVpZvpbR8gDLM1biPKopJRx0IduNdDX7PJCgSOEKlbtrHH5nPnTlW
1BNJzidt6skFfiFjfrEqKvjx1k2LLbUXv0S6zz8gGxPqvv4USZLsmUywl3Fi5TEPv11atIqxzvlH
UE9r+TJB6GTbcDTIqzCiAotP+6TlFSxNNsCUbjKvFZmsBdgjEESGHGHluop5VL/GnA1Kvud3J1k6
nwvVqPl2qKccOQsvJ7tQ0qvZksPzpFaKPv6EwlKX0VOivFv3FWoOrW3dbmWbwCjcLGX4I0+/mYDR
p+vLqHPlOwzgOPZ26FYOrvqE/kYUpaKul5Difm2sAorESRBWSFNDlTHl2UFg1qhnDhAjJe8au6Oz
HxLgN34vlXQa6Tn1xQsXr3m2IBgjccyYz5Umu3Zeq+LBcDZBN0KJTa81iEqVCCXr/S6NTBebg2DG
XQx/shjZr1JMMeIjwAycj4C+AsxPIC/mMbCITIpXpxIwBxI+4C+7WJrJpmVi5DLgo9C5y4YWaj+G
1nRcmQ3d5c75htQ87vL9bZLEclVFk3b/HMT2E522ZUjUzZQdt846T2YVIWZ24w0OUvZatLMXJKFJ
dBmAvFzn1JA+3MHv9aG2DBBR2rawPdWE1+vsgPQ17r2vN/DWtyt6DV+5G0v+LEuRQpeDi3EFjVJL
FA4aTJfeRdwvzNBQY0ERdX448j7abPZ1uo4n5pDh3NIVZ5/851pWckH75FtJZtGzO9qhnLWdIMtG
NTzelgLCeizOSj1bqJ2HX/XgZ/ww636nt8E3J5tupIY0j+Zk+8wCyyxMkOBMWCu8zXDZA3Jv88s8
kLcEEUIAP5OoE70MZUAMQ5tg061gYmctNUvl13vNh/PyBE14hKrWjvb2C/yyQMxJnRD22l6fcjNh
JZVYbFqsRCV9FwOzbOxooaHW9LFcG4Bxud7dsh0QEin3/A509vKMNW/+wO6eKIKkm16LnMr9QnsT
e8uK8VYnARxIZzWxtBut67nOQwetrMVUzxEfhJR3l8OiQBRPV1Bgl+V/GrBfoLAiBWdUDfLWeKtT
tZxBYZ2jPshi1M4vlAMJFCv65vyTXkND/oWChWmZBoCl1kL3TT2G6uzlb454UcxV2FDM2AmKEwOh
Oev5GhkPJjQdPWccT7r7yxkIPII5ySO64LK6toLnNQekG36gGrVzJPKGol/yJJbwMfbhikTzyYg1
4FioqRMbaDp/qC5oi8Z2kLwTSmZWdFHAGPI2JIybQhr1QQBikqTxdgaY46soHzL/xF0Ire6ZBmEG
uRIvWcfunOsley4PCF2hCPZUtoh2TJSP30F9A/x5XxxEujRjncnt6I/FBsnf+lFJCr+8bIUxbO8l
PTeJ+C5/OD6L4BHESdLcg5EVG4U70w9b4hLeRq02Ho2ARUQxEmM2alkTYzbXwUUh9Igqa5Bcgec0
qlzdx9lr/qx2dcvaNnq8/AjSSjSRCBSH4SRNsT6EEFOUKw2HAiqhvicGub3gt35Y4DC2zqDqf+ud
f+anxKqcHStIZoS7W527sU3OcP9lftsIOdeN5YZ5BfOm4SVTAMatsvEVDjL8u9AQ+G2pxoAwDVxY
LcAWKgE+iyh2a037Uu16q+VvIwI43qZCie37za7Nr82wkSpmHEgHXtRjalIlufsk9nEMIw59ZKil
c4KQCXNYOY9YjEr7m0k2JRIrVmDyff1YwXg2v4SVwaCmUYzfN+Q2+abg5foqEMKjSkX5io8VfA72
skpgaDxryempP1ROMfFHCvR5LElXPMI8bv7nic49RvFCDT8hwysjCyHt4YEC6sazXPWk8lElJ36e
p6ukgt9m4F1vfb3HgEYrnwSzj3JL+lTQRv0pGtSdHvrqjqIP87/GPvg8CL1lBgwZJu0JFs7Y5CHa
IY742yE976QGkdB6Aos95F7Aq9vmB01d7V56PpNrkZRu0sM+Ti+NFGDXInE+e8xq2a/Jwr5ssyy8
mIe8yQSSMQZx5kJ6HJ178ta8cCtgqPjmNIJuryWm+MikJpd47PHDbxPWicj+r+OWa5uJGtDR23fz
BokVAgh4aXUh2dTUx85MgSza5Q0G8egyDXMTVUT5OAvM3H9hTYm6FrISFvIHHugryOYOMw+F9T1j
9wSAZhi5dVn2gQlyuxDdwoBdHMXlflzw3pxMrHhqYUdvxjN2GIgCSZWF8Vevj2lqfazMJEZ+ujdg
m2wddkzVLKElS5/9GZa9WYVty7aeib6pDsO84EC7xwPn4HrBtBsGlRh7zjA4eeOXUVMfETBpTfle
DNmU56iWTQqKX2YIbVT9f5fpwnyeoJcsiX2CaS/R1b3SMMMyO/vI0Qa9mt0jBhvNL5fpeaHplFSr
aESHy7iRpYFH+uxiN+0cH5SSpK4OUjG69VJcWp8jTZezxOcsv0Dul+Is43WqCF1kj9MukgL2CwBM
s+pHfWLrRuBdtldbPPgjCGwuiERU95IxvN/SAMGY3DkKP5edqC1kZVoRgIPPJnOlT9kLHnRXxECn
q4uG+5hHJYVDysqtNZIY54lrU81CWkMiN+Np9WJG8ojJMERymQ5J9/UBc60ZQ6fD6D91eBuJwIV7
wQ1E5FwP96DFMQ0h8W25kJbxT81qFJSv4syltWW216CRDwdpfxGoZuUOLYlAtZOEbs0CJR63VON1
k/b+vxdjEVESL9zIuXPlhMXBVW7mrzOfRzrObACpbkXKMCiThQ/JTd+k1AJp5mql2mfkd/CPr6sm
CSiuzbdd9AKJxua+qf0A6zxoLZUaZVHKI8z9u2Ky6dXNgz/YFcN4ko75pPAFUsMcEEX7u/sqpqtj
HBzSm/Mo1nlW8h0k09t3zRVd0tVkX9KkmwhKIaM+69Y22K0XdA7SG2dya5PVTkpjVaVro0lEbl+s
m8dcpKFKsSOgTa4WCM3Yg/hmKk++XbUwckmGuW2ztxQLmRrIuBulrFI7waX+aqtdWxz6VvKuU5KL
tbKilFtXLly+FNxVdCcrX6spEE/GFJF67BD3a+75PX4TeIDfe0PTCXg8KAF3zbGu0kilFAzgHEa9
75MrZYLheM1A4iVXmw89hh1oPH7m2Qj8Jw3Nhq3ZvtQNUO45dIXAd8hhuzUTHXOt4L8tvqaI4p91
UGEl9uEJXiJzLtlJPLWYTCxZa46MAr66PfWZAzBT4R2+FTZslQLJvLDfpwZXoBfY9OcmW0+6CHkI
UpfqrGfr1nJBGfvhij3nfawcJqBI74+wOBe0h+L8pAEMGNJhWuEjEeUizLNVWksW6E1UPJwSg7Rt
3DT5k7FWr61cFVy8t16nKdAg1fIUOFP+TTwisXGHs4fQor5qUa7QAdxBqevPKXVT6za7pcW6qm7E
2ctXU+94paFk/RiBgbVaUcMm7NOQPUmZuWB9SN9kODHmTxyYQb0A0qluKLkFxfm6NnI46fYfrDUJ
6WMsKkA8IXeV9EBLrSipkSZ+tJ5xmVCjjAtqEN7TtfwyzICz76lB+q3//GnLB/Lt1Dbf3aIyBtId
GXKxmPdTQSHD8V8yGlydE/2lX4gil+i5YfNp3osJiiTntmpk3NlvFDzjiJs72+QZkIDwlkq2Ey0l
v9cOrXhINblAeuBCvJT4kBTm+q+5kDCPvHQgUAhDYOxMBmVpSd2z6cfpp0H1cg9icxWKCKNiLIfb
SNml4rlUdx29uyUj4ntJCee2ZlL38PQGo27wqhsE66NVJH011QXMWnl5z6XcTzrFRnxliT/TbvUT
aCwiQ/eDYgxyk2HJyJdkSDkL8fdKpP0ZWuGF/Vm7EkjXFudUtnI5vcIsC+x/Auq6QkHz3GkyLYot
1ZTQR8oEaQ3F7QO4AUSMe7Dxevhxd7ARy1/fIoB/izMeFCTwvJRT+c5qwBC82tu5mNKrPzqUZG3N
hIG+mYs/TegX+NKp9w4A+Pqu7ESbL/VYT6EnAqorgk+e2INLfqeNCQ5+4xgDbu/LMMmtgMY01UcT
THcTmQaIL5JCE1l/pNBj2zR4JFawXcLdR5wkKqCk8HW4B+0VOf1qgCEJLtnhpJYnhboTrXKgcJ11
NhsOUYbCLpkDZfjj/xkaXRwO1ddfWOWptN+KzZQBx6PdADQqHznZ5UKTlzWZIw6agpwM4Ieka8Rk
R3NAen5cCsEJfrPuxEiyZ2NXyxxbxdfl1jOB1i6AMg+lx9hLAZl4dvR4CJ0QRnkKDxfCSeITry4F
PY4tNfLTtreA55Qhf8ZxLKtDK++44m/gIP/fj4h9a2G4GgNvA1zEpGrw6nVsfr+Uco/OX6Lq2o+7
ZT5+FRglOlcwlECGx04vBBecuObPXZq2KQKXsF5fcCWyhmwpk8ciUiP8mJeX75D/ykZ5BIWZLWPk
BwmqCorLR6/wSJc6P7cai82MeLR1EKhJzyf8kU/jmGqonhNhY3rru6AkNlZsu3qLz6qmUQPf4TZ6
0HRPMSCLkQSm03dFTBOvdNBNlncHiGHBv/7geA8MSNpbmera/MZWxzgSi34u7NTKaa0Tx9Zd509y
yZTNi5ZzRqyWCKRwqcjrlc5VE3H86uNkJ6gjyJd3agIiuL6oRYp7C8+vdQ1FMUiYTqq9EJOg03LX
ifkpO0Ljy+8+vuCL1hvycT87+mmXYdupfV2jn+ZHLb+PD+m+8seKDyQ1RDCKEdIp6JFrlooJZP7s
+Ut2pHEvtMyodsJ88lTlCrKlAxj+iinqRcm47zVjvBdKmLJzersHyeTcelzPurYaVdYCzMwFVDFz
s63I458H2XF0ghKnEO6wU/Q4UIgfIgIxyn6E/CShybGNKIm+if9hYvA8nO0Gtt9fy5XBQq4gEFFp
edYoBVS7s7KK9NglAOeD1/Wa+R/CoBiwFP3n2Gz8eTPP5qKETPGt3tnE6ig3vZG/oqX/L9Lvu1aG
JlpSVCB9AOQjdbQ8Nsb3IQYUDmiyXCQGfEdsX4DSecZqTTr84ihLGAGU5JILY1qDG6N4SPdvs6Q6
nVerb48mZW++gMXKj0DjZKmKGp7Lxrq+JuqL5qbaEPJhj0vRKG8Wu81iy1JvFhigWOU7an33SKLK
cVlL0GfvoSMxS3vknyvpO1909FdANNsdC2OBgeX4Npfm0b8OqU9qgbjIS++vpWzGZUZBsdofgpdP
6PEyVqku59BDhfqpvsVHCguM4kjfXzj1QoZ5BfvHH3H4CPMlitWXGuGdP754jBHKlc1HSGrE3hRL
ahkpMJZYpLuRu0bnRYUSvel9xDQOsOx0OW1D+N5zHPvHvoRsucXRWV/UGoScrl2ykz7P4EfzSrfq
D5cGk5Yj73GUJibKRcuwGftl71vgJxw4dg3u/+XGHWbX+UA5P0pCl5wS5fm0dQngwH/GEPULuFDM
+47/erL0YGnni2qegz4VoKSV9/Q0VdctyNOyGwNP9r24IuyLtv/wsJgTZBOgmfBYNXFUrUpZfgki
Ks258Jn+T6xwog+fm+od4lUnDrA6rJsW29bzwC3qdRTUgN+9zWf5JR5RgmLI7Ppn3Iq1IrWU0pZ1
FJZt6I967/aJM9NO7nRukQukWkmxH0ZM1Of2ouQDpwmnORuw86WV75IDiymgEya4menmx9htX0xx
YVeyVLSc3nezoL/TV9WIFA12D1W3JDlcqbOI4XqjHYRGYVF7w1BlMTQof0SbyDwv6SrO2UnclNXN
tOoTkJop/bZUyfbd96JigvaVA6bUSq5VzFKWBUabSzFiuw4XpooWrMgLwhR79PfhVhYwx7IWFjSA
is0frTzeBYGBNXLD41ljMguBpd+dKfJZusrVm36sYFp7r3qp8Ge9i51xsUeuJdH9wV/CPs8cJc2x
Vhn5LbR1ypMjl1+XzrG/lb73O2egqIesKS0Ie5rw50lhgNlx1YxcIw8J2MzvwL4ahBD8Bq3Zuhck
bfwMpQMZHcq+ifap5gSaN9uei2gkx36WNRhC6hfcS3hQUhnEQWVCWjpgyvIo6g7hakhoZnEZfbkf
5Cxg/iUtS4PWWiAsku/z99dyEeP6QC0QIk1DRw2VVc5FG+VIa7SI5Ohpv0HatLXOVHZT4L37rplP
PKMjVBDV6dbxaG3wN5iZ4F1tCO6FYoOoZ/qZZuNseiw1I5NQqQMpPk1YEssnQ2YWHQPECxj6OM3R
HCgcSSRDwWw1kYbYZsNLuDiy8Oy6olN5RoUrLL7QmqggxNpiB8bPb7lhl7/wIfKhxlPCPB5wOqkO
eQKswE9HVXsMHDM2ztmStWpDShiBVCMAOdiOt3qlmOoSG89W9OQ/DswJ5g4Lzm4U/2lNpTmXk6LF
LtUNvngS9cxsejHI4eJdqIzbDJvihwj6eAHg6zZZdUepHYiVmK/BALFPhp3WMmdrI05KVErc54pR
rCbaHZlSzgf2QbUEPmqUG70NzW2iTSVgk4S4j16/jKJGgMsPSZ0N6a4jqzncuFCvc25jEJuMe/BY
rp25bk8bMbN0/ftvIAT4ZiF94KC3h8I0Db/L0iNuUOkPvJmi1VsN5uF0ARbWMkQuECq7pHY2ZJL8
MdMfgnWqybtmp+tiPi8vwGaO5rjlXdDAHnv0UDlQQW6LHQhoeo2PfR9taAf1lO0/CgUZA87y2Lo0
wWs4iD2VjP+hw8eldlbJIgfycmJCwkdJ4v6ccoEQiSJnn7DtrkLmGmLzp02KngQRgE9KRhKpw8Zu
7XGsIatwNPrS3RlCSumqIgs+Khn8cgxP0/MfHqVIHZHEiJy3Vo4UL8nyQ6U/PweCLP6AToe1OX+T
UkzfUOvQXKgRa1Jw+umAoK1pGTpRGwMihHwx1gifnwtHJa5yr6LXvU3igwpdNgzAqvO71t10X+Px
Jd8EVYgpnRKyxh+wCiQaYErtkDZDTRa8knGJv6NtXrI1+xA4LUPyu+demsQkNuviUQrtS2oCJb3E
PqZZxx+V42fNPpcHCl+CvFB4+90GKnLXGD82NCsw46ewmQjgDlr0U6glZMPov883NQWLa8yxI4Az
3zdY06G59cXQpVjPBKmfA57T8Yzzwr0l6K2qn/WFy8hyep9pEHCCJMIX5W7CBDkbuXuLZris67Yc
WCT2P/VG/+dgPcM+HXUqVtAZdRRdn0gbladT3muJR+vgtEp8UAr1XOi/v5lWLuUi/Qm71V9DU28Q
d2MhPF2uRO9srfY1dU7bXs/bSdpjROEDlembB2E6QyVDurY/opPfQuvfT2g2VWR8QRs905dRws1d
GBE6HD8BcKwqrZeLosVE/WJ2G2AzDEXjgxEP+UzeR5XdE8guSWjPSoNugaolmMFqbdI/DIdar2JE
zXcc2Ucm6Gc1DStTOIGfLg+Lp79vWIKnTG2tfFCUmNXPdnkb4orbAbvwVApLdH+g7yCBHK5xMKF6
nw5IISdGB0S7/R1otB2oBlnmVn935G4msHs1L3yn7b985tOq+h8KnndAW34icdGipOC5xIpp3gVH
Nnd50lz36SNztV5ueMQzXZD6xdXPJFAx3fY06ZvdSTURVeLEc2usxZ0YUwOA6mUMy5xXIxr2LYdR
e5CMV20efrO2WAsOPkUU/i5VmRJSWHrXRoP5+rHVlPikbfR4JxVGnW8Z7A/4P+lKt9Qhv8dn+hNR
UKs2uB5reqo27LXiAAvQVZB0L7K6uc9CYYcwJPSMTzdFuXYEk57VEAkZKcT5V+xDhhLK3CGBWSda
BxlAWyy4ibMAco9cFx/YEDFT450hz0newhy3CZc1ZAJ42qUqVsuCnTQoqSoZPuCaNJBiv3iqCJ70
vD3EIuB4XxWmXqhIeUaPmXfoXTEiCwMhMhUH90w5qbT1i3H9aYxEV82/ium24K3l1Rj8iWZKY78m
6nwu5XunC1nRTUKyp6uxoik1JPAqA0KAwRT1x/nqFQ85L9Jzj4pfWALCRiRckvH0078P0JkIPRr6
U36kt9wL6zuN5gfx8xdaf/4rAm3VMxVh6foYSACS5Fl6XV9yow53EnQ8Ft+Ugzw4mjrwZxLsnAhF
ovf9gcxn6ZYa9idLr/Jhm/c/SyhbFHYarKUg1iA4WE0mnsskpK2s85nWby6tvPYNARqjdYJGi9vh
GXpjYPwIaWQ+cymdbDtDbzHtFQG0PdWKaZuF0eOZdplU3YsgGLc1K502Ie/FtkRKn3UFjlA/DjVy
dXrn+1HaAHx4cE2K1dP/iCIz2wC1FLm9cD5V7O6fo/hH+Q5NNOYwdOEDmtdUenvYx5Kf/O1K+t3s
WHAUNP8mLv6kqWycqEWjGJqmU2rIlbz4OnGce8pDYU2RmH6qFFd+KbNakQ4XXudLDwuuuWECmf1w
2QdXCdtuuEHp2CUyfUMrEkdWOsbSdAlektTQBNdN1domp/lg73ui7PUWJXng0/PAzwJegOVbpOMi
tET4I8L3vulPj443DloVtsqTr+LcDhkH8bg8eUYDx+YuXyYzSEUdXFHD24wIRZi8ykzwBBtfiBmz
RWoaAFxFsYQ3lQJul2BNIAzKxYuYSRHu34FEhdwmClmy+ZIoGHN2Sk11fmg8lCM0Ov+YiFgdBNtV
J3AS6Kbe/jQYcO8dq7IB/EDLiA8anEbjdKsmNwnjRJGIjCLx6GxP9D1KcDQEZq6w2NpZK8Cvtpfz
2FkdP+RbaQAjdUQOUV67PcsOD3XwaE7KIqLebOl+M5m6kunaIho9thxiaFgJyuoIYPskpfC6iB+R
co6sHCIU2Ky8TLvyLDyTVm8JfgwT+2AU0thT3cN07TK8BRRW1TXVJ8NZFFfZUYZuz89wTKV41AH1
o3ZhN2kmThzwaZuP1z6rNiSakX1pOUGyrmY2hMMtFmFzS3J+pC2ZYVVV2TMNdLWBY71phEm/v6tT
BF3RHXOV2LupVkFw+RGt9VPUccUbLTVWGMvmGH8fwhvlfLs6zAaZut6+OcIQTZS/0DO4mv+2UOWi
kQgm86bwO9Xz0K3y+t4OCbKuMTq4KNB6iDn1rfGnNBeaxPp6eOJIvkQlUmSiH8GHcA+0GguZxpYh
Yk+rzuyc1eeq3XDWmvwP79hHdNa4UTcpZ0ksm7RgIY0vIBJDH1r3pFqJ2hQ9ajmOo+yHXUAlLdXg
IvTHi/L8VLrMvk7+64UZbv8BJ8Fo/YlLVYJ+dENg4xGzVRguJJbyETdJxCzxw9lgoR3lXYwGRQT7
O1lqc9t9hIPTr7DcCZYe5GKmsczew0f4l6b/LmwVBwS7i+i7Vw6jQUzvrGT5mNUA7sW/LzQQMUjG
SSr9qX27x9GpLdAR41lEB31QReqcz+UF/7Z5pdPiMYJYBWRHfUM7n6vftikXVj5PHsvvBg4ZtkrS
lR+S2AO4FN3QujiSShd+Uzo0KAWSCUIMz3N58SxDRwUVkSShVexb4xEB1+PcigB0YzFTuhejg2Bm
0LFFp6e5cZ+wVKF3NZE/AqfqlzFYxpxih/DQyn4/VZi1ieKbC7SLn38tvHSfWt6++mFbEODbDt1P
xI1MzPl7oOpdFHYyJzfcruoj7xmgXGVe8fHvoHSHXhG+yrEYWk5Yprbu1p1OTfAcuY1icKZAhebX
O7iR2enM6x2G2uKr3vogsnNOEcu5regApqCnsn4N8MXM16FbDVrho3qBZKznymmX8YlZQNlm9jqC
SbHdK8vpOzuwQQZOhWnwZxHsQ4SkqKNPB9WlslboVb86Zv2MiJOcSbocjweVLophkvkzD/fsEHfj
JNa5mTvLKwZTYJmuoruObW9BFkeJkW8GkWTZ/076vLZpf1MUro6cDUzTeHY91m8zDMlJ+dCBn78x
ir7VSEQDxDcaAj3J0KWMgra2OYBwydjosTQMcCeg/IFx1yluJDnpvnH7hd9qHUK/KznmjG29SYJ/
cDJ1YTy/u7xJitNETYmubt6RnSttcFuO+Ogcqw6IIfrDq7LZWuhruuxd+SwZFJvKVetUJsXMOFBn
19EMMvWq0AWulO2hjR+/ULo80MHRVRadQMg60m4ygxi8E9kl7g45Iwy0aFUfURBiUspiAnDo8YBb
EjX0rBWvLdxOo7czxgQtHbM3zkvi+CJWaMUm9GlQz1WIcjt68VVmNXo5tJbbSNJQ93yhgupm8QD9
JM/IAkWF1IxVOT6FL0xNqz1AWtuVQPC1vmgmfDusA9oF0ua7nDIASS4JybHuaMQk6E1KxAD2hPBV
RaIpoteiPZH+mHWDkdjF0OLVg6q2nSaH4mJ9lAPaWc87R8UmRz3X/fxQ2cgtUOlS+2IJPB3yQAkT
65z+zxnEuGgamreJq5GjKjG0pAlbuC6qYudn1Hf6Rxc1Thh08sT0k7eWlHXumV7hYfKQZeFiSEPU
ateBVW8zHOcetR4OsyuKiNP79hzR4G3jdNKWa0yV22yQJMyUsR2E3EwmazV3zzbHPbH3tJ32TShw
1vaw/R7sr2HzF6v7Bg/nuqH4ckFZp1jGB5ETuE0aFOA4kJlHNTof+6em9ZO46baDpenbg/4S6p1Y
jkfo97oSNbntcp+G4xLuKMCcB2I+WsVjxfghWsAXfrm393Ei4/F0mx8rmHgOofewjknrl922fKyl
fYMtx76nNt88Tl65QlI0nXjVxnqJ/hMCRKpDU85x9nZiJ6wqOtWHWHbzfdi0wCmchl7oWRb6f7ST
wgo95bhf+in1HKdfDUNRKfVY4LMvWThXedacIHeOZ5y87JZE+bkjse5hV5yio4eBuhOGkrFhg2SE
fk2UnP6cb5gOZJGy/M6bY3Ypl3Djy2f61bxEpxjBhUgqutP0JcolRK+GToMRc47GeWlOHEIOPY3L
8BXb9WpCc2pSCpxsEvf16rCBwuNM63N69i6n/hBQGiLJM2X4egQ1MxOFtlJ9oxTW9Vc1gl5ZvYru
lzidnc0Nvb79H8qoyJLk+lk/7bl84+Y/MCHzYwiqsQhfyf2qrVLAYfrtOfo/OuR/JA+135ADKToS
hyJllKm+nsL3rQH2NV5y+r6y9sQ/d3lBD2UzA4kwCPLiQvqgujfv/oVnVz0wMtHI7eyzC2/mKXu5
TIDASPHy4U9h/Nh79y8nH5jOW1FOE7PoJe5Oie0iL0HAVYOjvfhjePewjzDc26PDH94jZOm5JI3X
cAmFiBM+J2I2QfcgR4VOeqW+O/8v93Y3LsJWLHKRq+QrCty+e2JYk21c4o3ErYhc7d2bmEwhvfqm
xjp9NuzttWamee95z2d9nQ6SQFfR/0D3RH+A2t9ecgdqhzLufIvwLW2jTD/PoGdxp6N3RwAvcntw
BK6TNn/Ef9n862M9yIvHhTzwUygNsTuJNV1gtFIGcrl765QJ4nOe4vWDwyrct8kvQ4eB0ZP4kXwU
i9aMNs+rTmhbFwLexPt4hkqcXlohQoz1vhWQ4gw49CbWyKRrSuCnuaPCUnt2GeahD8UIlMgVHPfh
nYlXZe7tsSY9xKBv8xAXXhKhRNx7L6zQUGeYU+HV3s1IBTivs3pq24jIaGnuYgNdrZqsS3nV7F6D
C2mNUGirEJ4VoVU+Js6K1yEMui2MoREJiZ1lk51pp8RwPMkzi8sYsz4K+KXJ9kYNb0dXHYTZ2PEA
AycNSWt6Qnbp83aj2sQsWKD9Gp4XUMCpGIo3BE8zRZ0+l99ucW7jL1pkVNr40hvQnc0a4ApB3cVw
5XmhGGPJsXBkMhpchxhxi8fbaOzCSLRb2Yp7Oqhmv2NZjmy+MKfeu9BS0l4fVGBKF61efP2Mfkxd
qIghf9eLB12qzI9OCM5WqVGc0ed3t3fiXq7geB9kukgtUDH4npcDKNrqueb3sbIMUNA7OsSYvYEI
pvWOC9Tjjuz52Q5Gu+3Ip3UPS/g72q9pvyDIJfu110949s0xEXbMEJ42JWu1Af/BcU+BLNmzQReM
AzlvKMN/wMUYK4iYIHwVlJhqqpqzjUC41fdPV43I02Gs56Xs7E7egi397yyKmxV3jGI0lTXyTj3d
Hg1TSZ6JNpLvzn5pTNWcG8ysy6PjYYYNNPRZKM9Uh5grCcJ//CVpvDcyoKUGIX+e/cDV+DmVkybJ
W/nrSIIWR51HVS58QS4dT+LBkey1/6LwpUQwPJOh7+4zwLX+2eTS8XUoGjhKoowAFQcrhsa8zmSk
G3tNvJzpO7yRZsYJsPUCWOMvcqtU7XwQEFs3PS1XVABXGu+a9TIF6pqtuOe2xgFJKdt2cKbHT1yV
V+6J7dIKszGmmw8tfFZS6ZTFoTpoIToxcd1a/tMW7eUT0u+k35SbCjbqvAB1f/Gg6rBlFipfgtpV
J83uAE11BOvp52z3PplwdfpmX54JedWsB2NZAsdCLPbxRkgrOV+YwoMr2dv1Lkg6JQO1B4gP3mjF
3DO6Kvdr51DQXnZs4tzKvgNtTbTl9vmU5NdFrKxtwN/4Y+DSonwP9ju8FPqIvKBhHj4CccEQR2oi
lWKO+CmXXeUHAD+Up9NowlxMmypVnGLFKGUItAYsoDI7ckYNa2Z0GX1+mnceIXRj3kHmUVJ9W+DM
rs8WpM7NRbZY3N50kTTD0HT3AwaVwXm3SLgRbB2MUd6lli56vLLjOlqRfuJg5+/sLfoxlWA+fcqg
uFXy0x0a1uwyD3yJqH0KrBuE93GD0XnPxwzUqU9BLq0eH1/34hULesDVPDEhXLaX56Ueq7fJqVaW
IgCp3yMWApKIxbBJR3M6PJGKYcR9dGhy3mhySMCHpoQ+dGrdUbZi8sLPKHRcKiQ+O24HwtvXm35w
dlpT3VkM5arw1V/F9JqrXHv+Z+HbmAYCHF8/YJav0HKUvg6BATLNXedNE1iiL5/MZH0oVeZBMs88
/ECmbtHgMPEcgZkv+PL4ZSCNntAmdAdaTFBIgs7/iUclSzIBjZI01cwQ2vl3RzB9zmF0QLTuOZdN
s/ttBD9AQctPH1HDsJjqs7/35uckjc4jXat4q8ywx+HyPQMKiUb/ZS8AQ+cJq1gqewRr8jIxq2VG
3foZiLTJKcREIX0A28LJSscyTZlQKoWNuPgr9kStCnCpx9x5VybuHdaX55I2loEq0dNKVzIIiO+H
GZAUunE2S+xOJlF2q6ViLR4DEcdN7s+atFLGWMkeg6BR8+91vriAjTLCd9HGHgGO8LTK0EaCSNuH
0X3bbfB/An3Sl3YI6UK2IteN213GP0yokKFZONouIcHr2vgzTZV9bDCS+GL2TgagG1Or0F/iCD2p
xezP/Ra8nV7TQyiMBPqF/3pTl8y8cDUTW45s6X2sGg/heXijqC7QS27/DMO5SGuJ2WXSGahic8kb
zWbaRfbLPONAqoYdd+FNmWbzoPg/yIe/wdKPVspMgaaRI/h7BLiAWuR1KDGlVLfXhCRzDT1Zot/l
mLts9VZfc7esY57U5fx0wtX/0KSeCk2qMO+lfXzLQZ5+0m1P7jAIUyXm1FnSb8+Pngg1y4c8sxMD
/f0wsZw7PqaTB9D0dXk+g1P9VtiBZa825OzJw0H4x10MaZLyEOF8Zz+BymI5E4LKkTVtTzVdrhYc
dbZbkfxTMhhCz0TsgUfFuFKZLb968L0hfaStuLC3fD3yTERk8b8t5N6CIPSnZ0n6lLh2o8hlT97a
a3m+dCqmsdMie5A7dZ+uvnwK0LWUwIoCeYJfrDPZB5tNw57HE6SI3UF00fZgPbaYjJTKlBk1TYbr
IVDLBuWNUiLDTEKpBay4KYTitNjGCy5smk4dzMEnMOL4dlBaVN2B1xB+a4hIr73VhZxsfGUr6Mg2
NVset62fFPQyW4/89rt6CEy6iK0U/Y13MDYORiUl5w09x19ziJJiATUjgAPBNmBYZ9paAWTGVbMg
rL+49qi6Cta2pteH0M4qhErhTkWWeqKQFjad1cs+kCSxWaOwnkSmUDYt+4xxROSoEvFd54n1tUyX
/yiBK4vKyiNKoPLhITTKQM1Tqy8nwhBzxNG4IHwVL8iQjyhULB2KH/bDMrBhV7yHbUUChgTTHCDo
IRy31Zm44oqTA7jochSqrw2mdjThEvwxBX4iHTtDi62zNSLtFY+6fkXt0A2a+8NQbx+XRrX0HiGO
NnDa362WnNUq8ekUt7UEJRmoIQHKIUY3FA6aGQqUpjpsi7JuPV5nZaSw8CY0PHykX3C/IoddZSj3
xJ9tdxazm5thwDfhmeqz2Oby0kgMPPhdv84cbRmD7YBfODcsHYC1SBXP0wvFXpyCP6pKGsjz1Hjt
Vu2WFXkWCtmtmfJ/im9T0Ek7/qPHckSMJTYud78CEPzDsjz2QwTYkpZ5kZVHuTlk0vf4298nYyYF
ea9wTiYbRx5NCli9gje9Yp9p7tLbLc2iZruq3cpHCmJYXJQQaFwyfGb+B+31AQDjJh2E9KQ4jyS9
ZWzdtBq+YWZqxYytIAOynKL3Zv9phaTeXy1QpXlkxggiQHPXCwkgtVLc5CMNGWFEzb2kLFxThcS5
z9J2Ye9j4San5/4Ox+o4FrjzjttDjVqHRwACVn8OEAiOUr97mzb2h/c0F3Xxbhxf3zt8OBfkJydm
6Ah+jDC9lubpuIod5OWBvp8qsblwDIU6Rw+YgRK5DyJFZ3w5HFWVZWrbAaS91OfhLpEaqbGHxYLW
XNsGK1dlNX1gd5nb3GQUhvdNnVoEoMXxTsZ7fU/1Dw61GO74ljIU0GZQLkfUouhevv644ZQFFe0s
RIuU/mCsZ7udibNasKWhRcvGOc1UrQT/+W1gjweqS2Fu6X/EQ1NZ6/rYuAN+025PjzM25xYm4uZP
9YCoTqsZeBTET6EMFtc5DEjKrOh3kwqTIphgI4jnUZJkPQUYmv2WrIMEkWCLlQPCPfK1tjlg0slh
hDAJn9Ub46etk++ZN44Ayr8RE+A0Xd96+B31hya+DkOkE5/VNET1WQI3eF6ruo4bKikmReCnvPsa
fRVUeBujl8XkEqQCwYoyGLzYPyTeo/BWPXKB2/TYyRkipsXJzaQN/SbgM9JZfBoevymyXGo4ovv7
G3phxYu/+m/aEkbPiZ2RXZMTCf8aETsUHmXJbxmhlEbAsJjORvRBJLjwralhlYtWjhak8iFUMgWt
d+JFIds2JjdMPKa0buK0HjUgLEgslU4lkcmKqWoQxZajGANI209I/jrPYS9LHGu6nE7N5mXoSYD8
Y1NTL2Uf6UbKZduS3eCmQox8gN5LHquQ6nvaeJ+qKQBcV400te9FsnwBFndSbtz75OaP1AA96K0R
IQ4EzITpQhY6iha6mXPUp6mYh32HJl7oi+t8LM3LMj2hvVgH2qmHaeTQgTVBr1zbGj9KEnKx7fTK
jt9DYavAmXU0fdGvSMjI9RXciwxKDDKI1gevAJc4Wv0SjuXY3+zUojuw0skZrsrJNUs7M8V6xQbp
6FCT1InbpDGW43mygUee2Km66pS4Nv6fzu3fxnbryJY1j8nipzybEDdnEXUEdN/VjGTBYPD+IZws
gDAZz+HKioyxyhrONp2vfzpUTXo6DOyTr5SnTbUqDE4x7ZHeZITgr+7ntUqejZKytidii0h9Yq4Z
VdvsxDNEGrd+05g6jH7HAHo08LXpDRv0r7g1N20Wt3IFW1OsGw/9FkSLi2tBVwuBJ9ORvW+0G3OM
9PJ6nWf9UujnZkSdLHqkjaKHt3djvqDKcQxKufT5o9qDdkdOgocsPM53E6DUjq/QgK6XtC9r5/wb
cQZ5jew8g8Vkl1/R43+54/rWj51tKU+SEFduwiEU3Brr6VO39DMZH+Pzr58ogRGjSTsq+WWLfK51
PjyC6N2wj6JoFUPYsoZ2xcf228e/ga7+/SyjQXlryyWi+Ki28D0z8v9uxDnZtBaOnpPWuUleTI6H
AgrSfC4E0gH8tdWjUdxJF0IGOZB9u5xTo9LE3PhN+MObJ4zkXz4pEDu/aIMB6SPJFvoBZG8KeTvq
XIDqCPiz/bRzflTCULUdug6yMyOgXyAQl+HF8Z9l0DeoREuYUSdzp71vwoOPJHewbV6JSNAggZSO
bEysd2Sjr1CV1Z1BjC/OH4Wmypl7IHPm90wZH1Mghx+0xWH6vbXT4pQNeykajYKkwiXoe6G76zn3
oVh/+edaFbB+GtWo/o3f9NzVL/h9b49rxoJuKpZ9YqjIKMe+uQvN0yQtwO6xqpot358Scb+NhCTz
7hd5UwDN8gMqv22ldf2irnBR6gh42Y/KjpOGqHJU9S0UwWwLonXXR68NAeA1CWyIZ0Dddtm5oHcq
WBXsJVBwCT2tN0A7gQ3mAQ3FmecAJZGWlb2NMlEquAylGPtdqfwJLsel/YKEdY7n9VAdOcNu1hpj
67VWFDT50w5psWxPRUTqJEXpPANHpuEKbP/36DEFFk4XBsCyuWA9rHb+Mjg3O0lFaFtSXIOxrM+3
VlTe5es3ZSj2+CdgtsoLkTjERHHMtyfSR0X5mnzp1QzjKgA1JWdMz++Mwl86Qtzbj+35hmouj3XI
C+e3i/AjaQzwyi6bFO4k2ratqUWWbz1KUQh00b1bwzy5lF45oXaZyO5AgfgK3BlWVUrSD2RrSrLb
aqOfBQEwmXFuoYq8PD+Yqd352VEnDqcyiwDCAZdM177CI/SFwgJB4yX3XaU+BFHgDiTPBJ+5Vhhu
89rSe+IoTowiGF8Zimbf1Ko1qmDUC1BoJxGsFxVWGrXPl8UZT5PLB5KDGHaXX5Cfz+qYr8J2oW9c
wpkU6Kd8bSOpfNMnL9/hdk8Y2lFq3KEaa120EcxPhQr+R/BQ4g3TqWzVWOONZkBKVBN0gPnuz1tP
u+hGf94ZbwgxAdLniferLBt2HmvksZoGAde/roU2RRXxSMBenWdajAUtxpzunUV4pBEen+LlDvm1
oohnnA8WQG2casiX5jdodW2j7au4Lg5og2VEN6OmbwHHK4ISEnW+I7EV8v3cteD4J0PDBzAOiClk
DbR9SkCuzN7W9eDcRG8MD+f4i9VXPdtK3SZ/s8QSFFYkM4PKTK0nYsi64Og6uBuu8Mq6HFor6zoQ
bM27Ldl66Rruec1tktH3lYsGss0rTVukJ79UBvs7RluLlA74Ajokhuyhnh5SviqCRqKeyVayrSDn
gdfIHogIBqYnQzkwL2alR2geGYygKvmbELLXaFTUZMVuA88PZZUBGDoq9Ro8hSDKcehr5fis26m2
UfrGN1Crs7vOh8ZWKVJTHfPWE6R0WuDSM+om1DlTsSXLmxzrAX7Z8RuEG5FyBbbHfNVp6uW04lID
+LNUv6zxT2urYV+fDVJ/iOViAtywwBFG5f+Kbtddf5dy1QhQ6eCnmTULijJ5BD8eXaYb7+eqa3ge
GaDETm6T9Xq3xC1DDD9faQ5ZPeWSBeJ2QEK9uTVVJnAUiFTqhrMqimPoL7RefIPMXCZyddG4wPzw
Z7Ytk6RmA6wFWgW6ShMYYp+Xjmp9CFL6LhaTaAfBToz6+NBn2P8lzMhaVyPZI6VMaYooJQ9hOq8G
TqDYwbAFNw6ZLFRTz1tEo9JnKYcDLUU+RmlJgABTm9nY7Cit4EJ87/mAtxU5Ai+QzbVwyuSrvuf3
35haX7eMu1SvwYvboymko9lG3HxYj+eCHG/2ipkIqq7tN2Y+oqP/7yvSl2BA3b7+lhXaJtnT0aw3
QlZza6Pz4gYHljba7nTVO7moOTjKxJlyQvbC64jYi6YvbQAozv9yhyWe+ij4pYGS7cOGKK85Awfr
8o2FHobwBbQjC//rFUkIoSbeRAbhmYJfTzYXI4UHItDWcGvjsGdvN0WGpC6oKqua9wEaLvyrwGvk
LyNMG3+0BAf+V7hJhbD8h5i4LGcIrPzTI/ZdBR6EbkpFnEiAJELOo//qKLFs2h3ZU7c4e0yKf2Bn
vMNs0UX753dN9iiBj6R5VCY1mu9rsdbboRfGGqAfJ2aV2M8+yhdxjUgZDuO5T6ZXj42SfDO2AJnI
F77qGjtIPkLqM2f0ZEqhefi3ea9Mfb+IoryXXlCvSJI//6w0XEdlN/emN3luqV5ZYxr4PtkYXw6+
ffhgSGXd4Swsnd48/mTqoMjxxUW27YGtlgSHDBKMP2eR8VE0KLvOlYElatFW9hMoViw9Sh5yaZJN
be19lO1p65BMEJvqb2UXuLoX2/OQQnU9R8Kjfwrj8mKsqZITz3wEAXua7Ew0+bd0Nvu/OZfmCKY2
Jug2o5XqiSpd5C7pE3ymdj4l5yVQUTGmTFiKo07SQqM4jlPYakJtF0GEPnAD3YWcOSby6ODR3Npq
bo7rRHLTMImadkCFJeYJkTHYAXl7i0ioi/5yM54T1QrLyw+Mozp0E0bCbCdTtR2F71ITKuKxwpLT
IEVq/Gp35hbd3vzYfeFtPtl537aziW1LPCL23I3o1LfWQC4asT3bVDiMaOM9g6mFS+gDENxJxaY6
h3iiUpHThjIKb1IaDfdWsVYbsP21SLIlCLV5Y0Df/34g3qKmY8grkYs4tXiF+D8doFpaduGH08Im
WJbCjVcdyst2tk1ASZveEa/8v1EmUG9bVVL7VN76icedWyUuswayoBm7iwRxXuSfmLxcBEUOUjdI
xMHVnwSRHCRYVzeOPrmfBZZvGXCy6CeE4fcaJgPZHuzTC7wZFLJcjyOMtYfRZmZ6hzroox9lWav9
ymnRTZ96v3Z7hEgL3wPffTdvCZrq/JZF21KWNOWb22GSpULe9b5C+7UGE9stDoezEuSsbOasmFI0
jYCdvTTwihl7f8BwL02C5IMTiwsGJktJBB4385KindalLusCtuXV5G+FbjnjNho9+Zkd7MWy7oyR
kS5DzovoHYicGxIhzCjszy+jQV2XjvNTaGQh5zitaxY5+xQY/g09A4fS+8eHKtKiWYYH9qQfOBu8
T5eOAsJHyhBRA6FIJHX5Sqn6PAKvUdfaE0lcUmnZ+vzjM8R3Vr0iWTGJGsF6ewPa7p0Av6cZgNIs
uoB2KO7vo9e9Xs7Whcz/hgjFwJAIU0HY4Clia//0ed9+JsCTzdY0z401LsMurTnUKIy2hjUu00qU
3ZHza6e+8z/VSy8Nnhmnjp+ivtB1ZC37uZlqA3qqsupHLvsioZniyugGDG09cu/wCEIK1C/RIEJd
LAOPkJlBLUEOSfAAUyxCjo7kmDFPp3RnlzuOCwKtPM8+Uz3xsX6/Z+0IGep2o2XjKfyq14wirzt0
ydBN7yP5ZXE7B/TIX1VYFXFE+7D5aBwmgH8cZsq4w75e9euYInAf28Tn6yyEtq4E5lESnWi6kefs
OYODc/LkQakDlRvGdYbccf2r+HvrtqGq7NiCpcd1jNVSVAPR/245tgIAb+h5YdrihVfb1+zpKgVj
j9h/7yKgtzXgZXav9WkD/embCbiRi3JN652dlGweZ4t7YLv62nNCG3fOMoyISYdKSZIo1lZi3e/S
15FegF0u9jVk1dHoGxwQGGLhU4oeZcb+cdiDbL+gbEvMe7rQmz5LXjDY3qo+QNYyXc3eEY7GFDIE
oudti1okrYpAPm3j4qMlVEUVlpO7chYpeH5DQcrSlCDsCfezpzVIreNxZ8C4FeQa8y2schp6mnPa
mqQa7jih2wFjAM1KUrh8jquH4m+prNwjeDAdolCB/nsvfC6/aynaJDqz04lKMSZfaDQx/sSV0/Ao
gcfWCEjZw/jF4qEiwXquc6v0gk31HqTzXEsR1DKbg4VNhelHFLjv6JsSvlDHT7LgjuqQm+e4PCwx
YSr2T84heie/dTwRZ+J/0DbBb59h/QBPTMJa1it/465e8VYtA+v4Z7u+O/FoY3ExIPs89A9coZhs
KkgL7jhzlGEoTFgxfgwgo0asgZu1w43Hf/8DVP08+NWjRlW4owMoohv/XpRwskcRkqan9gPUIUDL
8QGJTGiPaPkKDVYUBp8iT86hkq/YUzuUNZMqkA1+RGiuFJK21SSE7uPJurEDyF6toXyAODQpPngR
WbplXMK9Ejslhu3oqn9rasNPlH4Hl/umWzHGL+R3Ob4Yd2ioemVmhSVaxdHv3bUMYCRxEpr+SG+o
CYjGM57YKFZ7/K1MQmpL5RFY/1ZURppR6ifBRv0+g0yRk+6lycnCvR2MWv1P6SvSC2VlI7Bgq9A4
ldmXQK57BFOUECFH41H7Y92h2gzXl57kcA99EQ7Ac1bqWHUGFxdr7YeBo235SHdYSoOFGj/Z3/Fv
x9quvyHFRnJTyOudQx42705HLSBq1suBVsLBdfU5EpCHrGppju+G6EeoS6vCVzNtIds/Un8A3Zgf
FwSja90YsXfQdeDQo5Olb91kvGb4qfO2OlfAKP+wK99gg4fgRYGBtmQ5WezN80eAmY8rY4Hf1Xf/
xZjLtQrUExNX3yaoSlUTyo23Rt7sSzp346CBEGgFGTF35zZNQylomm8MgbvPm/6InDnbWHR0Y9o+
x3UXO1JSDVx3lLIkdDn+jcQv6mArA6ua3TJbT8Tf1hpBz/zTUUQ62e8Djr2YVd7YEMOXWkVYl+mI
xGhxyaLro83OktHgkWV6lkBT6IGms3yzog4MUcf5U3NEtcbhKvRm+xyG9yzJjvvVaBxufT4vGJUF
nUNCLm2j892nWaMFoGCMBIwwsqy2z7PzdVyfDKklMHzdxxx+PH5EKmtNTBBQZ5rzML7XR6GkxhaT
Y761/+T6nTpTw7BSfYCJTpeklyEu96KD7UREWJRSy7KaDVKuhhK+I8k4Gd/K/cCaHfWCcpRkuWGe
kqjfICTpQkeuDp9tCQCDmFb64E6aCbR3zz2P2qLjLI4Ov35ADuAFYZvrQ8yz8c9n6rgYWiXGzW05
7pFrb9eTL7HeZIhZuhbmAXF63gM3HehEhdrERyJ2XOcnHfDuTNF3p3abq9YaJLa55nJ7/0RfWWNp
lRidAdIgobnvyvNjH7nUVDTu9spfUPHthgurI5z4icya/sxv2ycCT1rgCGEPc1lsdx1Cik7kZCHl
pJpvrT+jrIH1WMiyQNIC58n1tuy8/omeftFe64UCvC3GLKPoDmcI6iXAZptKTVbXq9m9tS/AUsV+
pkmGDkfGW7JjaeKwxzZ1swahadjrKpoOP8oE1cgiX2ndJHxA59CvQI0WD9vx+x/isFibvNRllPQ8
IjkKW9S8p5mk0dJyKoHFd4nfUQ2t68qcJhPU8TSrWy9aMKMIyYRe8crvj8KIIsmhDelBhB0nh4mD
E4et4w8g0JuAdaDmLBuUncX/vkoU1siszATD0CLZB+IOSB5qpfAMD20/1hOLeKvkCIrS+tqnBLQp
oV3Ctxm+z1/v72RBtRxf8FElirdbQf059gRNfpg+pA83roZyB/pfWB7Fx18f2e5KZpqDa1hgUHQc
Xn4ri9JrHzZ8W0UomFhqYon1u42GKeiu76+f4/uCNAN2Yq11ziDFFAQddzgJTEPdf4qvhdUj5JVi
yKmGmJ4qfX0T43AN8aLVsXIVXUX3qkF7fHCMsmxeiWVfPduA4Ym0r1WrdbrlAm9CrNLc2P7N+Je6
YJQq9TXVDW82aDobrwWKL9dw3LWQ0Xbb4IGa02FG8Grk+MhSiUFJ4ui4dAxYsgSpzNJ5ZwDH02T2
410OR1KJdryRUq/Zdo4TZhU8BL+2jZZ/dMYgVXIbjJ9nXLnLRgli0suOajH992bnGT7eAmoXTf5V
/iC43Sd3eerDbcNW0x4QeNF87xCk0PZhfUEdzpcOGLJDbGXbm3E9PhP2ixErbzSLVd+B75yYvK1d
nmwhrZJsnDdswIAfo9p8nEc+HnTkeyOQI8pE/rDJODzjNvS9uNLdKkZjXAS+zGpO9pX6mYccDK3u
sGWR2AaOis+MZcCYXm3DNO2FLTJEVSjYIKHhgiNPNNDiqeKtkM8djUt/H+k5zLFRac/8Fp4WbT/G
8j3aj6GIvkyGS9KD/QS0uml8ICcoSvuAaqx8pLdeLKCVdWs9AsJMFq73/PmInB6ZKOrAYsAyk/iA
+mKE7PVkuAHIe1Z4J4pwG3zdiHZDRkPrtLswD+M/pFbHVkN7M+UAh8hhnBAO+jNFFEKdABnHcG0r
L/OoVAt931qvaS7ZWXQ6i8hYNaun6wExQ9LBTwbPlYp2JTzoEjzTqR6VE29IBa859oLd64Obfw9U
Vd+ro6xO8l6xAN0c+A/tFM8VpBZOjuO0FnaifdpZ29xzKBqkwAxIQ01Ndo8UPjekX7rpWgWQDTOY
ghZxBCKozfXKDsFF0RLjwFOEDkXaSX8YQA2qRy85vPJt6XkB2DLfD+eoBLMszSsmpx8+PclsEJ8C
g2Mjvl97hezZjigVqTq2/69G5vhfEWVJ+brDrZqo3qUaxT0GrgNichfI2bsm//O0/zsXItzY2rZf
Lf/oieFd+6UYyozyrsVb7TdZm19Z5p4Ykzaaw02xy7rQ7iZbWxrk4oQA18TKfSsiKf0F+xnD0vrn
xWXOoe3tElzyRv0URaNlnhptLogjlSo19pSzchvdO3RVo4qdvPQUvENLZAzgygbHKQAb/P6DkQbY
SU7z3Gp7MH/Q42NBh7REIQTzu6+poqbfnWITFXZgBJ9xGyLH+ZTsV1dJ7RwB3YygrS6E7naQAjue
/dNu/iHRN2TPfTe+2aFku3XzzFeTLdvIMlREzSEJvYGSU7f4g0A8FP29SER0J8Ow8HrkYJF3xkK0
CZFEE/FY5EsF0dLOS4YBrCd7FZF8Oou9dWGe5AhPek2mNP/wyPaQxr580RTzeWPrtP7R1K73AKEw
3tNQHT54d2FTZ9V5jOePefpLkmQzapkySMu1fUGrlVcqsEIGpoq9QPEI8tyeQNXMyJw4UedEqEPp
uqkUOjQI0KGmCUK5Rrbg3zUL2JSmaMfQ8i9JhkKH/mM26/tRH+IFRg9m8EUP2R8kUd11jGTOON7I
6QgvBJGAwD79/6XGJLetiVJQwg2C/K9rzTDmQjUEw6FO4tznmGMh9kN/0mXnlvQu5GMo8NckZ135
ZUobf2QijMOlmCXfD2iy8YVcJhmEOz7Qh433zi6iswN6r7l/pDNXfFTVc4bZiLZwfqUV6362HF13
bPN3ngU9OHN1gJDXPoToQUO7+1UwUFfv+6XiE9xrWNO6XdWG5s/Okx+uX9Z3OaRKzzldPPQFcDow
YoF4X9UryLpVwBlF3Sl6GnN+TUZLD5yq1l80k6YMIqku/55bKPyeWKhALxgVEre10URwY9pfMuRI
ttXlWboE0Va3MK993Z7vkNLT4FmsF9pHrLhwKZ38jAMm+63Z8i3o5GiKQc2Z8Utm3c6deooihMFr
AW0ZeoHaflkBwR9g8I8anGb8seK8kwy1UfGSj3qcyO3r/PDuQAPzRr2ZXDdclsUBW4XQeGyRKjYM
vRMFJeCrtkCyszMJCpItbVXIwKoVNsM7FMAQ19bezmzNSoBw2gw9o3StCsJ/uZHmP1zdj8HFJyjE
okX4DVl/3Pv9RnIp414rKmAxMh/X4bp4AHAXP5Ttdwa31eIGLpH0T3hboEEIY0C0CE/I3epZJBzP
8urYloFp2swt/TbHDvSHnSP6or9bNOjacchvbYHrSUYooh5bulmih0oKPnoXZgYF5nbyFT/cdg0T
iPI3Cg6f7MgoE1XPp8Vor9epHbKKeptzEkjdkMwXnLdakoymv8IMAOYjVnOl84cPFdC7L02oLyPV
Y81F88u1URbQt98ZHZ/N8kzNhGB+TrAaDbdKdP71EpMoost59Y0bmVeNjbOthbDoPX9ZdS62T1MC
URoMNGm0XyaonGtI692Zo48+LxbxZNskQCxXb0h89IqeOW+b6OsuX33sexPl+WcPQ/ItRCAj3pu+
MPP+qRhUjNL5q/ysd70kAaSCzN0b95gQpltrFQ9/PFhU/T3QS+4kB+HHtgGUgauTRDJ+vk/ls9wN
ua9aJw1IxU0RT44YsA0zuWUgaEh1ZUhheYQVO8sGFUgbE5tn5iEyOZUKPex14+5Ol/czB3NotV7M
587ifkIy9jTolPAMQKnIuF45eRhjbdsXpPrlg1DyDA8JieDonMAb5XYIbVc024+IAHRPfEJrR76L
Xp/UEEy1WcfBGpoVPOKZDYXOqQW8bGKVBoGxfPbX/G1QBTuzlbL5VI93m6HSMhKpWYafzpN4ZVWI
VR71vuQ32oZj3cet1Oqg8ySmuKm6c1XK21NfHEReflm1BK3eQ1psC3joUQHDkZpUcw389Gg4D9rD
xN3o1TZ6hiWSxXPkerKywqwpkxtoruQsdw/Ns4tCEjuUK+Do3R4qqce3M4Yh7pqlpq4Jfbiax+fE
kfem2w4G1EBSoUsaKXd0Ye3640PxSU0gOyOXDa5AxkSRjlMgJqVhdlfMF1DsBiGfWMDotQze8h/a
ptoDO9bL8sDHn+JFMvBIXUljatySK7WulpgWXxmFsJRpeZPsjUNfknrksj5TqjbDcVvhoXUP5fow
1RgqE2lY++IWA1mJkUDUSlrB2mRT2GbFUtS3DVWKxu63v3SXWDg4D5RCeVrqNBE7T013m+wHHG+B
DKptf9/s1wz/djVm2YJsHjwBTHlE0eA5l/xwdlKVFWraa7mq4ZurN/FkeYkrzdUVrPD5h1Vge18B
J9kI6mUjAaAsq/VnugIzfnIkyeqjyKioxj6gWLI2ZDbZnLEQcZetJNn2m7a7heJa4S9ESStD0Jz8
5ActWC63ievgu1/tBmQX3yfpoq3hwzFm6KN3lHyGONFubAtQKDndoBQe4usSjlR+C0WwQAjUdOB8
Uyx7FR21jBRXRJ2JimJsQu3Wrc/qIYCiuRqP8jFVN6BB6BMRFhUoWyr6rLKFb+xgKh/cuPM6gOvB
RQlccDYPrYqI628Vz0ZKGcltcgEPnT0IVKof4nPIfC5wW3uQ1X8ky0Ie5Ed+yn45q41eXbjST78R
HZ+YA0NBgHTGqpWflZeXTOm7f2O2SA3webOOmy6bhGrs/kZUooVWWLtvzzrVugJDetT44bmrWT1b
t7nJpqwYDMWWpa5Oiu69fMsnpd5Tht9xKPGRUi09/9Md21rTYX8sTy7luhbBSKR1tWTg85IDvmBh
DPTG9tT370pdySZ1j9z19yEkKCK2ONmxhKuw+yUzX1LTlzZoMtRarJX3kSWman3EbLLuLslA8cr1
SrQLmhaQqg49dJIbAJOv75p4HEk4pvbyh8xSlk5/wqkAsGw/YJYhT748CQL6dORNnN5sErqDRH5O
ZgOhX2g1xrcV3bKAp5mnfeANi0QuUKT6hjIsPNVNREH0WFkc9qv7op+m0CGde6S+zKRhrvVncLjf
DkdYJhZ4s/hAaB2nkP5Ee3iP9ilPxiswQFMbq8SqFfueOYOMMm7X55nO0MKpnmc9V+qZojpFha3d
LR0pjZMq2454KUVUMY44J87yHIbpHZ1yekPGKI3BT57qmo9/4aGLv16BEa7LG5B6xnAAymYYlunE
nFM+80CG/7dzUhZ9PQ7ZxcvUuPPlEo8BSsvFF5q4SFwpIIZWZSQHERIvIaGRr8jt0Px0zkc+ywfk
gdsVcoZLmxWkz4uJAeOhgafhT4dgD2WgSZI7gQMEkN0APHbRXp2K+EU1r04T2Q+eG0eqlers511h
PAgjPS5XymS8wGyjDp2gmqH8tEFCFfgb1UQ+j82/9Gfb25uj4CdQ8TelOfE/PGHOGUjdNbRIggqv
dra56PzCGztr8kWzpiTDgZ6VJbHP8/PL2jGhchVTFuBMB1JqToV+vizkjSGMwfXxdMYa1SXPaDza
vxWAeBsJJAmSN7hpTRiYVxFLBqz0ypMLlpUKOHdY5QzOL1oYI2mmklnP4iL27/rW8QjT3zA0pPai
Ulg020aEwaQ8+RKhdHGfY2cs/xKXxgLQ+4nLc14nEmxMTlO2A8UObz9qun4JzxO3YW43CmuPRx54
27NRYDIol9TCxFN2lTQmbBjGSe8Tlh30B6J0wi51K+mHnBYEi+xfW/d8PTjDwjc2J4G+jtpesa7T
5v0YBa1PGJHCS1Pzm05gPA/S656F1VKKdXCLc/AMTl9ABLo+A9whG6Ap33LiG6vs0LvyemcOJ2SW
5e1jFV0v3if8JeTENeobdfkQ0sX8+DFdI34peZosGK3cHM1XXujF4DY8/RakC4Rnxfj5AVQBFwwP
ZdinO2vgaJ4JCot9pzPbA3h4FfncBMRACntCri22ytiHyjph1scJSPXIGLvjYYokXtMxq7eeVlLd
grthVa//IBOkxiR4PJ+G4mSKma7rT0ZKpfqxavG5PNtKrbg84uokQxlrcBOv3+E8GkhdRT3+1tLm
10/SvcibZeNeznnNhqkgvrhfd/yg4SsaK+fCKn45oAVxxMfkcEPshoEeG9KrGG3iIeORDbryUb5p
X4sFjYkNNHw2RGRGSkL1yJnuZiisMAO9zf4dDpJWR/kgy/fNTuCLCik2bapEH65UoP2RGlaFx3hl
xjgGeNja66aFktViquih6CFxR17QB0UsEm6iCoTBvsm5tNI9vn+Go5NEUInAuwe34CmabKKFxMpU
87Kg983w+liT4X8AW3RNPyRUtlGaqmpCvxWG52nf50L5Jnwb4uaVGuYH6c2vnYaoF6dhZs9B1X9j
BSvGf1HmCXSC32ssKeGodSYJBqTZEpO2GPO5Fv3yfrHkwu4Y/L8Abrn3ld2QOOwIdmErH+acQtLe
m0HL+tzl+ViRq7e9yNoJKwXRVCeWS1DhXWWLIGPkMWHj8yNtB/S4lMg0XjNIFSzLZ5NvOFrfcIPz
mJZwC9yuO2gm/A5x9JYzsUdyaru4ISyOE/Slm0N/bvL7ywNbM+Ls99JhzWEDaausTjiP5KFsFX+i
q5mJrvOdafUPzSzO2GlV2Dk8CUQv/t+xNLAONIY37HzX6vStXld5T747cj2zWlxKr55/oQ/iSwSe
xb+9Z3UYtIxddApP2rTcuPwOLoLs6qW7WrCOnLAKgmjBnkAU5OYPJHEfGWe4xPSYNzZcmftEsBJq
AmZf7swbGQ2JbLnNmYsEoOl2nWJduzKAonhlCR2Jv+DCcO7c//sgdTLUacgK3XvdzXEEFSwQ/7tP
vNfAY62dg2BvGvmINJJt+YylTSI5ryifQz97Wus3DWmHs0La4OKrjXEV1LFsTuJUQTSPqdbJckD7
m8C9ii8hSiYa2UiXESsLR8hy7n9BgimYVtHJ9PtltCw1R4l+cCc+ZU/v3jx8S8BH99fzE6d9ThQQ
XTxFIef7Py4r221/VxJZXFrJHWmjY4T9sgt19Q2Ge9sNkIQtzZ+bUeviH4TmhclX4u9woDKH5BAl
xNSFmQ/n9TTE4e/s5ACedXcyKjp9j0k7pHoxcB8yDFZcx7EUblHkiNqhIojG0yedxzhoJPz/enPO
4hQ4jz+uzLFCrDsIKjTHNF3JcQNro7TOwbRiBGxhz11AJGLDI3zS1sAoCnsd07ZhHpFsvsi6ZhYc
i7eJMPkJ4/WmUp6aaEo/tzwNgod+7BpxQMZhuUqIQYaOPEAHMKHNOwoH+QNm5CBPj5fTvOFjZOGI
AZ80Bb0FLdnc5NV886kmi2nSdKYWs5smNcHVkgnGZ6UgpUO6KRZxof5+XVusMUSSvmKrj8MqcuwS
7sna+6EU4/TWcyIaXAVXi4/sXDagLmSsWtIQ7O66K/uvu2nut+60X48azIood3AQeusDagGgvKKS
VT0MeN4zaYjNYtjzEUARVHRis85S/pX+OVlyU0Uxk12Go4zOlvZfA78eSQilm+5IRTQAoWNzvv+g
Cx/Uf+uaAhnLNwPo80MlCilVGoHpJR7AjVw8pw4f46qxDpy17V2X0e3Wci6HVNhddmM5a6gOZT4g
dLj2MEYfbEnoMlEP7iOtsjm00ac0fIP07xSDUd6qLpy/gTVMWNsR7gZVsv84t5+Qw/EUvLFyQgXX
2ScL4NY8EQkjAXBUeD9b4yItG6j+jw5AZct8ga2z88QVdge978ZMxFwmNwxoVGeCtrN3So7zZtVj
Jq4Dhn8a87fOuzLMAAvKlXkZZghv1vuhoAtbqUDC/NgXF6NpDhFxf76fg1NN3KGglJy6f6aRhEXv
4SaS/7U4Q90lwiTzKds1eUZkW9yH8AO9i5JeMcvf01uwshwAPRRSf1ZGrz3O9vm4RwAH6uSxq5ln
GlRlcCZcU3USlpEeB6s6AL3t3AKQvdGafjMK7nj5Sbw4IKeXl7veuBT4Z7toseOffihPpApHiglg
CB4cIg1YJXEe/9ioiCxx1yDSqj8WeaccKXLtqWEaq/nkjehlvtZ8Sbi9BfmYiylOiMtM+b+yb5Q2
NjfXmMRJ1DEmAs8qHrfvCknYe22uzoGkJsORqZxyHdDbK3ovIkR0T7FrV4wnKqoAZzwMp3qIh+Qb
oeIg1mcs8hB3nnvuGVoe6bervAK+TtDfxwJM6TXmGPWUC/L5/huoIhu7DsSZbhm3dujlh+4Hjxfs
+VjiUTJGKCx+ugmUbUEgdyDwEXkedeyWEEo7SfsPE99AFBw0jIX6nz5LWh6hgZbMlzqO18yPNZQU
KSnm8X5RtobRy0a82cUGoBEKWvyfuqM5cHORN1SI2Tl1B3KUGWSaKbEtt157axMT3WGwIz/Ya/4g
ZuJEn4lusQ9pOjOw6H3HJUKcZtiCwjkTwsQYLTxuGUink4Ymcn8YUR4CrRoWQVbpG0c6B3trzuLZ
YigyPdzOgsY/66szymsyS+/xSgUFuTW8cqzMq6YnjyldLZ+e/0C6/QW3Q6bIZqoWF7QM+lx38mMU
fYipBLdSydOhLXQ2P6Son0z0mBKGjRtI+Ds/Xbht/pwiDYuzylo3wZyF0AD3Id/hq4oTbyPqUQR2
t5jqgdpqrkikgnCIvztIfFKOF1plR6cGHdx35KfPKiu1y+NY4C+OaDtLiA9gYAr1/lgCiFQKfien
nQnChd2TeGtwXnOT5vbjIeSxOwHwyx0DrbX5vWjBCCXDlgIipQM0a3fDJLj5UdUtL+qUxKhXtjge
jpN333Bo2KveOaoDs1+ek1FHQBdJ25gYJEw00ONjHQ3ghpM6TOc9FysDDFYHao2bz6ev6z87e937
WyGrAIYTDsOK7GrFDM8WuOjXgPuETH033t1ZaGwRbWF1y3k/G6G2U6U738pL9JjJKggzYVqGJp90
JWBPpy/LsIhxM/3UTb691Z4jubvv1WDckvd74VJVbMoePQPtYbGUa23EGU4S1KCgZ6yYiD57KXpK
jWORJcC6XgdkrGJ49e8Tm/sHiYtUqtOZWCO6SVhNLJY8bmI7ZYigeZXYo/d2hI7xTlTnninvdXz+
4x+MfpZZbh6UUHFIfI5pkpHUPTYrT83MPXCnp/UAW9yzvFj2Z1TIFf50MJAjdm0Dcokx1kt4enWi
8ghSpgEcS5z9uiQlCrC73DkR6zhSXwGi//zAmEQutVeVRSLM+v9YtFC4DkZjjS0BrzdYwvevP05S
G6cCMx1RFfyzZdMqujlbejua5IWRYnbVO1Egou95cBZZWV2wPN9kMx8xWtUrzMr7JVlG1Nn6E0D3
VlPfQx17jeqgPgPl/4cHRwIqw+3PVPMZtbmibMFstLEeU4gnbxIv5+8n0VBfQs+giB9Xj6OqiAhC
C1ydTbo+CXI3R9p1JEY8ub1GL1Atpzt2o7ddUdVaEGxQV9/eMUnzms4vHX0dcpT6J4mx7fHGxdqf
v6nBC0r2SEOU2CI+h5FGdI0GQuYna4uVQcXwxXalQrECInSdt5wC7xq9yj0yFj/o/O1OsZhgsd9n
w2agr63n2DS1ojBSu6oesQ164T939PITrATJCyxlQZlwR55vnsYqk4pV6Gn9uzORJ6Ucs78rUM7N
Mdq7AvG6V7R3o3dMrH2yGRGBt/7TtdCHhl0qOQ1LLg4ciU16FO4PDHRo4G/RuxCutFsMl4jDIUor
JHQ0HwbW41FPuHqcSfFpC5x+W5AuDI42i8g8clihkIIz5HMZ/xS2eLcNMS2EKREveV0/U9iT2wTN
6vpynKNlO00KN62ffmWyr4w/djOD1aEyBQRPvUJ3H1xtcglKKVPWOWl653aQYFfn2Amrv8q80MTi
5VSVZr/KFZfk9CdR+qgS7HKm1mkiiCSOAEjw5MsJuGldZ2NLxAfKpwPBJgdy99t9+cjo36k0iIik
wDWHBBl01kE4yg6mWl8G8eJlY+6wlqVmS5+qhHK7RVJuYLZDTIlkwI1Css1PjjGM2oGVSua97vcC
sQxvBaQFw6KH20+VrjGdETZoC+z/WsJ8Y9xQnzZLXNvpk/yGq6a09cRfwIyKIYI0shVFRZgGhhNp
TOoym657thp6uH0spSDHfPvEFNz8hy+CCf89qpXuygK2qjNdSR0qu+EZwEtFvWzTZgLu46jiYIWo
sb4KYvIlhYtF1t42X8H+zSI4tZYfDwz8Pd+4ZdjwMt9UanjdAPV/HLXJXg/k5woSMSAQUf14u730
ZvfBLV4VfqHKkMAMBxItZibfPBpGCz8A9sQMhTW0ztF8c8jmFKcPxoz6umXfeHHVzMSvFotnAzt3
Eyosx96S1aVzrdfhcDATewxAIFCHMxb4yuAXHBXhFm/fbzimna4RGdBfsd4nOIqqj93jl+XBc4EY
pOBubnwxL1RwrPPABoQa0tKx4x4NYUBU0pIE1PuV7rvfMm86bMGDaLTRIOQcfFGRkadRn9cTtaYo
S0eqHsm50LRgLmKPQAb+xklxvTVL0oAt5zh4pQC6Q3SSobSaOYLwHQTIllriLmJAora9umGpp3qZ
fjmai8O1/yZ6wRiABaxyPN3hZAWa5ijU9Pb7lYeHp/0XIe2RdBqW8jXSUb5QVNEoUvE+xCI58x2i
w8n5ejQNyvaDOUhsW+XrIwlacH9dlIWJrst4Tf+xxyMQl34JYmkJQMC5STKity8tJ9Va0j3/hqGm
3tpJef9Xr+1mKqcIubi//Zc30XJp/CyAH2uiQFyGVY8QA5KxsONyxpKVBDEiN2whDp4fRrI0OFC8
28Px7ajweVLYMspnpJ3PYg3lXEp2XHHigJnuSneBnG0rRRy6dFRtbI8b9oy5it4uADa7nEHRsfsT
jf9UMGsZYEY5PclaB/jZJOB4yvsk/wohp67hgdDI7ynysQXEZGu6V9guinVBjVMbHtVg61rgM9c2
0df+FNhjUNgUhj5YSho3C5EvR5mEbSv7GK5bIe8rX6+lXRRV5N5JvoBxkO3jrsQwd6oYK2Ddn2Yd
CKFdCQfmqJRbYub6hAFLLqhqWjB9Y1pmIqD6QzhPper4LNsTUHm2Mn+1Yu30RuR5VB6nrlXskSiW
v2GtF8VroMUcS+nuax8gYYUCZNSPa2lUJL0eu9K0hic0/kctSrTfsq2JXu0qQ/VLy8wvugFUkCqo
aQrKsQ8hooj43UH96hble3BgzygZxLEzjBhbz6HDUTvQbRkriwLntU1/NrKWhu13qQeEtSC5Bp1u
gGrva2+l0HQuhMj0CFSeW4E/f0yXMkXth18RX/Ez6R6NtCXm+fpoHJQTLIG/dY/R8jpgjXiFeVhU
QsZaodP7ICWW///RjcFSiIk2/znyQ/LGTXdsolcumnYxU0p43ngIjgedm8Txed90e2OSWrftpnTr
OF2ovXqzS7ep/KbcWRiaVVrJAZNKcjiCfSKBbxu6YlIl9TKdsCmubC30LdC7GiOqc5RhU0k7T5BM
AHKtLL7Fo/tGUvPhL/U/MPZC/QqkDWydLXAbjWjgtK36cWHg+DjyUzeWnTOil7ZFb8weGCgWa0gW
LKHxRlX49iDZ0S15HXUqzFjXqotoF5vyB7eSWYMY3TjEEoY9WoWxxNXQtRsGe+dcSUPpIDd0CkCj
Aj5IFuUefmFfqmsUCMFIJyIG7LVz2bVQIVTCDLMl6VmjvRWn62CmfM3EGP7ntDVEenXy7L3fpcIk
6TByH3IjeLyG1JfS7jVBLfey4khJs9U/+zlGUTaPP+rlXyU6yTdyYYccpmw95ZEGgQB6E1U3K/E9
0gmtPt2gNTFcL3hu5raw2GFUhS5sjdeYHZY3SwlJyuJwWkVmIUWIz1gLQr/3jrM93h7vd0ch6CHr
2r9iq3jQ3kx74ABXLRtPSWbQLhDFC0/g4NcJEmeQ3AkygqQ7MMzNlOfbi5kf9ZMRionT1/1ePXfA
FMjKKW7hABU/PXiWnHDjIVwX+eRxMl4Uaqa1xuyZk7XKpi4Lz3ycdA632f4dLjrbGuRrw65zemeC
V+yGhPPot3tRisWK3H+L4vkCv4FcLDleric0rbox1xsDL6WXXN3ruHR0UDvyVxfSaAPw+JFOhWi2
7T4l4nuOA7LCBqcS048/AMzqlm7SN9yuSK8StDl2hjMWT/OHYLxifr9mqWK8TVhwRm4v1EqVAzBb
Vz5LkuvX8AoNwgcfnz1yflTpnhYBPMTFY3YqHfBFC+wkIr9jFSgBbR4ErrAOXanCiuYTFcIMXSU5
h/CLE9sHEeRpjRRePmlVML2vCEfc46EtUJ3tpgS5+xMD+dAxYK+aJuazBkM9W6raMBpN6CyRiKjI
k1jJerQppOeQectogy0Ab5AMm5f7JKoVxq7Xo3cIXM/82+W2MbhB784bdTlCW2gcytxDJd0smZ5y
imqVVcEErwQ4UUF1bVx7J1RZg8pvGkVXm6SgZKMQ6fYFcXWGQkI6YCfUyH+5HdknGDwXeok0DOOZ
ijuVa01GTqwl5i/86wFW82V35hOfn94NpVGKrh6biLAQq1F5zrDYaobg1XJY50OilAbdWa2AJ/Aw
KEEY5WcqdeBB01Btu7swh1ntMR63QwHmCAXZ5aagDMkc5EcxdH8rxnA9rbY4PNpJ8bB5Ezj8EhmH
PCOw5iC9B5D/3zP1kwGqpb2igeOK0E7AnjkQ1lxR4Nmlb1C1qfIMK+vEiBiBNsw9lcqcUsmZxdOb
X5RkEI+J+o/UoLfbxkYLe/qhGI2O0GH18DFrSIMpX8NLIZirgJetq7lDvlAa+fmJO9E290RLi6P+
/eGS796nGY0h+UlopDug1LSkIuNOoci2VBgc2I9z6XnAWmZ2UaKtAFkQoAwzq0GBFRuw82MhIXH3
ob2Mk+NcTJBBJQMfVGNVsgJM1rcsNuUM/ecgkY9HvbJ7WtFxZaqfMzColYdRxQvr7NLQv1ctwJ28
9XOtAdHdpTdVVogljINFrYxT915gkhjU1ctvySv3d0joc783DpOKwlw4VeqHp8fP7BH+FMeoE1mQ
SU7UcaFMWmA2StIIwWtCQTv7K5/3kD8/yXT22IVp3QuGSzPDQAUkR1e1kasKB/v/Lf7ms8j2aTlU
GIJjz/B8wfk7NIAk4QPFnvTsuwD2jftwcAsgBfdTi+4MmIT3QAyVSBHJnWfP2EK2/3aMG8PUf6cS
2f84hP8b7/tsvwz8Oy54aB30oL2hrUgQE7q2tnXwGfb+o3zS72u0Scihx5Vqdq18hcDoVMoFZ2W4
2NUurFZXmGlMDqVD2mJI3TcABqon5Oovf39A6xloyjtGPWYvgrxSIuEzcdU8FNcvWuiPWgv7EBGC
4tloFcyhB8eXQX9aVbh0BXWy0yIbyUokNohj8iNeXgDvfykMSE3yBRwhpReeB4h/lKpL8+LMd4AS
DQBJCAXCohGPvJ6xhfB4RH8lbqgBTPIy4WtU53GAyloAA7kHiw0Hn22xa/wkl5P3XpVuCCtJEHZ5
+Sb6lklRpnpYNlx8IMnYIuQgORlSAH0mb8VMG9MbNarmq/pERZH5EsTD5jYA1h18OBzOm1tJnT3C
dXh4Z3ftO6YFhy2bo5hmzJpwAOJF7e2FeapjWOWMtBAIOzpMs1RN2xSOHOuZTDu1KeNxbg0KJryx
HGhDcQ2cAKZaj0t8dnaIPICkY0qjAWG4p0iyafC6E1Z1BXHLSV5K1tDpiWMtjSvAgwE9jtMsxnHc
WwEaEAhB3cos8nDR7owyfhjGDzFkUl2dvjDPtBWcphLvp23dOoR71UBPAJvLLKBkx4h0aS7NrY/f
l4Xoe1udVgCSHC+V+xV9MAKtBnSUETMv9k1Q05GCtp1kln9LMxIaqCbsvmeacx5weg/IDN+gRsvr
m2brlvE2YupqVDLF3B5TxNvOXhbrq3f5PHFKed1BpCEJivdUMmww8QPMhhjjbq31sYFKF7tH8fv8
EFHuk7r0DGakZ4nGiUDnjW+xG3V0B6j8+LeojsKY9BD6PR4wORY+jiTnSDrNlg0nkVWY5fXRsMxq
na7Mh2WDMBZLk7FQZZx59mOHDUhxhcJmngXw2/vbBaFWvzaKGbFVBv+jg4QGfnyFm17mt74Y7NW7
LkX8oY7sCauzB2gWofYv9lEkAi+WF8aQPwom/6CviHcg4a7lx9bWAA3f9LxnG85QLPlk3it3m6NE
c8/ZCzebMga13tZYNY5i3kqhELfAPY9kIdKYdQOLiY85ABOgAPUIBxpVFTu1me1Uv/Triug68v2M
lNvD+Q5GUXhQu/Tvd7KgA9S7D0mQUgX/ZLDvehxZ96Dukins/7dRTq61RmEMcPBCpmmDPoOcAM18
etJSbQq7PrD8GgwdiqINCNbpqccEd9/6fN9x/oGiQj2Fb+EDwHrhv86eLb+ZPmt5VgpX7txvDSEg
+0hZM6rncCjJ5d+grW69/P2YRIxzIryiiwe3bmPqRdNoaUaaGoaLxvHToYAfvBuQNwP2kgSKweCu
3eFHDSdb46eoO+CAQZNtDzpaz048Tnw8xvjhoCoau2W+YdOfnGn804EyT6yx/t58wAmQFIIqk7ig
kOUnL+jp8HQoWpi/AABE0zrw967EC0ipIt/QNIFiIrd/izrjzXDvMci7EMITdq4y9HXrZQG/+AyG
ew8eyZ/FXgZ02fBqb2DKS1SVWVr3UIuroctf3bma+7YbVOTBlxobmG1315ZD0ltuNa3Rynlv5Eiv
SuOiaoXjtEneeiUwy2DhVrZC+6LqPn8tgz5VLEEbIkfANojy4luHUhjtBWEq/H5+IRff1wGF5bpX
HOW9i2TPlp+63ZoihV2QMJ0XcjZ5ew25uUXCVKLo7ucKMGai5VBDgfIBSdfZA3zeDbP7pzZOuXpI
MGK5fIBQtB1YAkMUyifrE8/9jfm6IQ9ZYrhzxV6f5gKFV3amcbkNxIJxvesvswG7aAu9JbPrvrUh
3Eq53ECoymQlGhRWVl7mVGzEsprAq8VNKFDN7DJxc7m2/R8Mg9YFZGKTxfvVyUzyQzf0Dv+s9pF1
lk2N+ZI0Uj+UoMptPChXCbVcS3jJfzMPNUdMhSgawwE7Moid3gU9esRc4/zhcf6aw+3O7CXT3F8u
54gnWEjT7lT7hjKzD0Gr2qLNQ1sVckUZabVS7zJlOEPZktk5EZQeqHr8+IPSCCdBW3NxWOjwom0e
JhWlGVg7rRfOsuu7ir5wXGIMVyDQ06c8ds8yvfH24OfxXhUDAZMUAXYN3WhtmjY8U4usXaNSSONZ
7NrjLlp/AzL2siBNaxo+4C94JV10LJL1iNr+JjLAP9MMmrUcG3DMiw65Rr6L5KXVVFJTBjXoQ90E
fTcV4ytzxnSsiGAmnawWTda3J73plUGLebxlurZ41LERUPfkmWPzSiOkMcoI4XNYcdgWyhJr18GB
M0xmlJb/FKvtGoglm9G+d9VD4iyb/cpv8C2u/UOFZGJVLdRxhEzZyka6nY+7APmLdCC0tCbjkDky
65G5+598Q4y/xyONPNstPjzrJ7B0nG5hFUmTnVv2aQ1lbROvtxdLtrfOIOVWGSsvrj/th9924jtX
+rrcDbzkFvGzIUZpd55oL6MW7yWlF7LtbRc7Y2TMDSUxvG/uVa3LxD0yxF+UgsP7SEOhJwIWzmki
Ffs+o8u3dm4AYbTT3HWh7KQw6zcvEJSwtGirsLN/+fqH3dl84KGMjRRT5OwGFek8VQlbCtvoMX0F
jwYAqdjYFbwvuewybl60a2pRsDLvoWqJxUlnkYA6XkvK63m4h3eSjou7AV3vQJuX3eJCC5ih7FxG
EByhNIFSP4ozpKNFyRSQaUlmmqpYcvhIsYQjxwaFbYK5P0AlTl3Jzcp0rn6hfFRO2M2jCH87dqMF
NABue/aZsdTAJ+tXvDrbjnUTd4lKFTE1Vq9NHUQxkRw4mEevkeyMnYjHj2ZAsySCvZAtCkE7xURa
dOE1gpmXFVCzriKakYAj7Vrlndp8Z7RKXji4i1y8eF075ZV632/Xx8mnl2Dv1uN8DtmNV7b3sQoo
Xr12tfHoeuwFrtyCpLeHg66fGvTxqSv9M2dpCLNumoK9ahBoJaAU+8BeMTQZEnwwda2d26LxNNOL
IbbYDvLER2lKFD588UAQgQB0B1Riw2NGZDgkuhtMHlBYIllpcb6lwR0tJuMyuG8sPITzf1RVmePR
ky2xDsraD64/De1ICPzimrVU25OXp7OzydWSdYFO/8rs9jFzjavbap8273sfoV6uvMXs5PALfDMw
SZEAQ/6yCREtkgAfOyu6i1728H7IgtfLOWB6ahVeTNEdqotbPYZSuEYuwFAtJa/IgN5B3lJjAuKr
6Xd9DWwemMSY53JtFmUq/TY6zC6CIFYzpnTaCSY2GQuufn+hKBFWU/Py+huYpF20OOdxCXuYeTA3
F9g0y/kXA5BD8z8bZnBaoC/MKNjxQ5g+UEBpCq5XL2mL4/qm4tfIao29YnC0oCAE4ebyu8LjFDeq
7vCplK6kcMD7XAoUXRdJwr8Pe1N7ZxreNjm3QwrjVNXKpdr0bvbx5cdDr0K1AKtuEOmqUHwqjfl1
3jUytfZ272yWgEmC07Gp+7ij5PvbvxN2/bn5lZWP3vhEKfUhvlpuiyBbU1ye8zAuJEFx+XSLiXR7
fsEdDDTTtBP+o2YGpUM8/z3Y0gzdlhh9meunVqYdcUmgxaOUhcqF6oW1QUe5OZ3gySw6VvHr+xfm
48C654ABhJCrfwAwfG88ue65TaT6xwt4OhWA3Ybxiuvp2AkpSNVBGo4ecEkTPNNjsajOksZfdZ9I
HM8WRmRHE6Et1wxg6xSnxHxwVFyMjU2HMkICValGoGa1V26/gJRsCX30KNto6JzfAEbxqbvcSkYE
ON7T0dGLowzt/fMGPEDro1vUMiN4LbY/JtQSRWZdA1LogPvFuXOZoVo9HWQ4JW+Dv+LYouF8qdYD
NysFPx9X4Esa5sDqwL7K6t++uLkgaeqAfUw8FkNLPfxwdmEyepZR+ysGI0S+B4MZA7PnNfECM/jQ
qyfZVjSvVZuI3kTj8HhRkmwJt/jwCUlAKDtebKAP6PyES0BVCnhpxq7aCEtVvPGpGHEhEhDw368M
z6Uqb9XhgV68gNOHHsfnAPm32nXBtuFNZNSjeL0UJQi991OU/Ay1YBk9dCxz1lKP+MskJVWBiCCL
rnX7W8D3TrvPOOKCDNvCR8Irq/mqOleYPw7ZY35Xbb+themLa8bcQcq0a8ta9ehAx1lbaburVcv9
zWGC/+MSpXnK962Cz8o9mfWkJt9hat9A49EpOOQU9uPWnmkHcrDyf6cIIvS9IsUvbxjGD+2a7+Pj
h1NJQq89R7/8QYFA9xlfwvaeemJkF+hFMjL5MdQWotiyx6jVH6Y94uiJYDsWpazINY7F552PImR7
4J50ojnthbrWA8dwchG4HL4yk7whHaXWDtwHwozg8KI4OJZcpG4FktsNslLkldK8BeDZY8cbJm/U
PAoJ3by9cPWq1a7Q9T852O0DQf6eWPfD2Bcm1DDZN88qhxDWlBUw5bChnrIrGmmTu9iTrHZ+3EFX
1nLroZZY5O6TPlFoxiG9vvCXBGhyGWXBtqmowKlvZFNx7g/AV18jfKXb+g2l0Y172syLVtUYH0AY
fpoy3+L0e19rJ2Er+ZSfHf/qSTf7Z3QCXgJNhmiOQtvNAF43b3MbwKViZR97si6MWHz/ohiR62ZG
sE6gjK4KKNNAG2n2FJ+XGn08MKfTcsRX/j5knxAFJReAamOfNFn+v0HCmeYdjkpFedjQJZL+8zcI
nN83QlAqIJ1vsY5rHJUTXod9oMwbW3WG07VIiE8cIx55w5WeD8zmZjMPPoy2/eDMHsX0QOk0oGEv
9CIB+LLdC8jcVBQ24bdg3W7gDB70aQMDsWSvw4LS0mDeNhqYmuYEv0EINodzmPyrSeqwnNG0fbkF
+Annl5OetTbBsYS0wVs4vMZ4joNVo0CqvwZt3f0wLYY23HECKaVqKy9ndXeIcvpuO+u8ZmxZkB4K
zHt+fC6JtppVWiecZXC+/Dr7UDlCEpPfcRWHgkcq57o13w6FE+iQhXkMLhTNYvV5GANsX3dn3vvi
XortHgAeMCCLDxfUUv8XMuUVLpJz1yVj2JUk5xRYCZE7rM9eYlxBj//VHosJB7euLe7ROW8eoRch
0TimweR90vaRFxqIpS7gJDDTvOGUAyWncAFyJlJvwUI+ZVCze9uIgHDojbVtUnjhnX93dJ9lhAo7
4lQ9KvlVYXmM8wMLGUCi+dmTV1xJc8+raJxtziBAXbJa6K2k9J5oprInkvdoIUxXfy1yFLql0oLO
djA8YijNoQ4B+BZY1SWNz785ECsBYEFD9CrV4KayU/zl6fmpw3MvCZbXcMlkvex0y4QAge4/GcOB
rk5MUJNtpjfYD/xxrIrb0+VE86YeWFa2il+RXDQfhHlmEUl0acWRYE9lqGzX+TUmUgZGOeJFi3M5
F7rDZg8nNDS9OXB5v/MeWoV5FGe7DCQTDTUTy2uyP4vi3silLHOzL1Y3rgfQRr72KHCMc6lDdz9x
ocU6Zogtk1VDlSRw/v5Q4BBO4+cO2xeNUBoBoz6oGCZlTw+cPnCUeNzSlOMT5VkGrL9zOFwPNKf1
cIAA3EFtXpXQHxAjDudSN2OJkFs7cZuZW2f8Fg6MQQg4HvbAzbD/jPQqwN/k18ASil2gWrP2kJnl
/L5nrxyZKIKFThQbKd05HgLx2iDpnVc/v+9P2AyPXN6VORoF9NbwBWDK3hrv1A73/RnfZvECIKub
rrwYnmQJ+lUiuiIoNeUoKTjqnmVg24AJPLSSG5e7TwUY/QLy0zg5IA8X3yww74cfMfWGyaoiduxd
fa5L/L0mvAsUYIJWodVksGXCMTy2K09WRub4IzGfPEMaOxZn5ZcO2gngMSsqfuvuwLtKUO3BRPYc
e3PTgg9oNLrtYAO+jhtZjrhGaHC3ccSkHePnV8f8GsZQy2ifgwR/Oi1gz7m8Zz0DSjwSQEpcuTFy
Duh5ywxIwfdSv1fGN1jgy5vSAY+uxGsNYFE6MwF+ovo1ijdVJwkxZohGTuSp6tu8TbKoXHKA/+55
O9gPymcLSEYl5JCJIo3h8KQ/YXOPVbUTkKpZ0nmF0A4YOrt/eTt9PUhQ7jHuirH8SznNul5xrpbH
hF7KeXfkFvAC50opH4Ag4pbD4kwcz1P6wPwZwV94ukzJz52/csZSxOx99sLdwUmWLcVoWIIcTVAZ
8b3GiL+vnd3IHDoa388QP5ZBX8xL/pmhPMBW4uJjfrnAj8EdkgxDgFd1vf7KKjp3eAWtIVY2Xmtn
RPeevVH42B2bIOU7AsF/a81J8tO0/4MCuebNXG0XpGdOu7jS8TFol3stTh26IZCO7In8MC963hgB
Dq5uvjXjI0icK6wJ2V2piRGkJJ8HYFSWtIl3yQCsj00EWkYGW4r2bqg8KX5RhFIB+L7DhwajRrHw
/YgrMSDlffZpqiK5G75C+zBFmflPmf/DP6H2OZzVeE6dC/gCHOheQZI/lKU3xkG3i+BKitSYq2nU
yybVV54l1VqUVdF8Ct4/Ds3OSuE2Lontvi0ognwYOGDMYdR44bjvKXtcAWyqVrw1mz+JKqEheoTM
UJiLxeQtBQc4eD2V6bIbvxyw1yBRA5jWjO+ypJ+YljSKxLNxbdkuaxrApSLRbEWdbtcZB7DTU644
nuGy2I7jyWLxbUbD7ovYQ+vOn3q1ngahv3svBVcpzwiy+DUh4gHJ8pWR7DEu2jjnvQGBLycOhCXU
0B/6oiP4rnwlHXPNRGxxgtFkGW5HcHctz1fXIqonu7elfN78Ov+zHz3qaO3mrjBQf0TMR3bcUcuK
PE+ArN42WbkWcKvrUojCp/9loxqfKs4Vwt8ffjmUVlZLbmrvFow/N9aSv/csL4ru/ZXf09QhMXAf
yeh3ysikRAj7Mvc2cij4372eqSng1/SuYGJ8OTHDmjfY2sGi1wybGmvQXiL2ez17n31AmrTadBcs
ocVyV5VFSvS553nRZQcQpcWq25GKuqLXo+fAOKhtJ+xTFfd/N6Z1rDTsSI42Vn9QccPrEdy3VWEQ
1b2B63UsIpNGnuT7J+dmFpS78rAsFXn0/00bKfpZmfPYyQRe/9G81vZbZy8gQxDUSZjKnRGctYkU
ngVPjly5mHGNlweKK8UMPkDzfXQJ04HWaT6+VduHd9/jG34EDEAUW49OkXdakewA97F3R8Tc34Qv
+y+LT9rwapun2j1uZlPKadZK4Bq3H/05Hv5h17rN3MHyILZciJ3QaaIKBqzBQNLczw81soOyy48E
IaS5N5OE3K4wLj/yUWP/r2Ajb98tkhgUZ/iuaHRrb8hz/Iy4spIRmUVLiuXVAaQbrwg430IwQoEv
QkhXM4UDmyCauliYrWwVVuxQtgdr6f3Bcs8Nx35f/l7O/J5RnkpXNuWKwRuAapB5ccTft045qyOi
y6DV/t8F5okK/rkTOOlAGqqTl6VawzY8yrehf6ecbVn9dP91dwI/kGq+sFCzHJN880mzyPPZMTYB
5D7Udl4rhk/TigA/wBMIfDXBmvT+Le8njHEofSWexCZ/W9cGDnjrOg7g+LeoMQXBuRwWschUZKF9
EGh3o+zZA3zwmXTVojRiPyxVHCwPHsOKulMoBrqPb1IV0JZ4ezt5kJX+tQeeqn7Ej05dBkz7fWHt
ItiDz9sNcB1kxFWvhKwPxhS7ec66vkKa/8cuXISmmAtjrFOTCTi1TJ/vzuCNXczz7f5zBeezBuGW
13ZmJJ1fUjdcrb88BUrPtdGKZ4CF1Nf2oxxdXHMmi7tmFRDsFVlK7JMIBohXaKrxEGc0emReNzTk
QO1MmwSpFafh3xKJgF5GoVipG6yYBYSV6uN3v+HQug8pBMoFLiIB7rCtyT99uyTlA5UHzKWC4aP7
zsfmKyUUHMbCYbSDqaDwF7vlNEyonDcHKSQnpiBxoHchMCZxcpU/gBK9pB1k00/0t4FMiu6aP7Pd
3USEv3ON3k9TkutzTI1zHYSyRAmgC6HnO8Bb+yaWaBNE5yjmdNYQfaHLbdMkf+RYPOXMRPGp587A
0oWl7mNTltZWMcfnTet7bnHjgtnRT6D1qsq1t0QZVcOokmUqKSheQvhlfrpKnGwk237hUPhEu8By
9USQBeZuhygJ4OCxptxTq/GMIYgABeR3gDhU8sVDfsOMHms1M4dCSNrEB+tW6QuT1/skS+ur2qap
oLJeR01EFkE5gtp8Ab+N45Y7VUeB89ai6GTX3uY94Y1+c1OJBnUsw5QYEXWH+hqGUNTkT9fEUxnc
JabeRvW/GACaJZ3lb5b92r5RpHL1XE2N6U+CgptNWKZnMB5U8uvPLhmmN+OoOcNiHityGNTOe6iA
8ZtUfLviGXNRImV8s+OXDXyBk3ieFxk1UlqZ3s0miL8z0E6DU/W3IayWb4gDiC4hRKISwTV0yOZb
FtesNbAHLgQ6IFezBwmSGbkAZx2PpdyRMbfIS63Kbu3eVR97FFWLHr4AoM/x1/d1PQM6CG09umAp
BVqqZ1hFTXYIOKsy/jtyInkj8niETBleFT6PEBHjKKMxaTHyAZrv9VRut1xvTPc5QrXQECJZg1Sg
hl5qSN8QPNInIFqJebfpK9zCiyG+jgNQlFVTxorRO9NWAECzpv9p3tuRPQpTkNw6DgcFp64bCzvm
a9edu13NrdjxfjvkMBggkFXkquIeA4IAIlwejVNB2FWXKHJvdyovuyUv971+On/Om3t2CFqylLhn
3z4BS5Qj0be2gYfxnwrAxLTVx0P4RJS9fYWxSrmaTbgZEi5+tTPB/We1wxxoMs/bhl/zc2P3f1Yf
e+hU6mBnWmvuwyHrvUfVypfwiS/6nY88MNbTJo5y3OBHYMWgTy0OjqTolDVAv6gqj/EPthVK5YKz
BaG2gyr2AkTZnW9AYdTQABNrWXqCjmwa6lPkKN5Y7uuHLKopDXF8bue1W3YlruMzWJesjfYZlhRq
pfdGIk1WUut4r+PmN9BAjE8j+IsdDiHVSapdNMely02Du6HQbl1uK2/vaPFTNYC5jnmbfO5pWJaS
exW8xhRkRZm+VSLMQELN57fa2D76wGAf74TZ7tViMxMTHHcumq3YHXC2eOwUycdtLUvrBRRgLCTD
wWrOgkKRzWDlNU5Hsl7hmD4opY7+KasxHKGrhJEMh/9DL2A/1kr8JwIagaS1peHpgeKSxL85UdAf
o3ZmL8h+ATqUggJYgS7uq0i+riqofDNCJJLhROwAF/gUH1sCclkMXnl946hA1E+6unQtfULa7Ask
+A8/KJ2FiLXVCyJdxx3PzUS46A68xGUvb7yK8Ztz50rNCmwj5MFlPIkUR4wHpzqQ4aBOCZ4Afz8E
NoND+JWFMzbp4By9jyqZCudXApCYMacqfab0pDZy7rmHyJJTawWF9McVcUxQVYhKwo5Ci8OvC2oV
a69YlZBLruXQNWfOqCdafY9qbbPR6SX1JVSdI4ZO0wE5d5/qfWXntXAi4Onkp1WcW4JcZmZPqQ5B
JD5yO3Hdudr4sEcXzqwZfdYi3rKAt3dW8z36Q6roXoiHfhJFlb3/xql3AdM6wgWE0ULmN27jgXeU
jZaVyZQfVl+znKnf5VgbzgyvQZhQp6YmwuugSO9iEAnwTnoUO1I+rTXF3Jt1jLMIPEFnn0jAn8Oh
PXoEHeqNzKMElP+BKvJdyefi46TEK3tLf0yX/oktD62pA1/B+Elo/7iafHggvIChDt0+7pNCeRWZ
sPdY9XjQtC0Tn5Hdlh2dDPjMlDTlpvt8Uxb/VFiOtbMNWWphHO6QyLGWnLqpsyUkZSekvzVk9I/H
gfEbpA1dQ3rdUS/tQqxr2vQ1bABtwNIVaQPYLLBfxjCSJrRM2WR6btY/cMPtamYvU9TnrVE9tn4f
SdlEKA0pPII2l+rkFm32J/emS8GvkcqWOr10hw9ouvt8gH+TI6hDCRqIWKJYOcpV7A+8/OR97bLx
Y94kpYHQNzfxRrUgNkfYZCnSi6flZ85PtjHpOu7odN+JVFE+1rGK7863fTeZLcurJi45zHOwG8YG
SvI6Dsw8ihAZNeZTC8DFDoV9GznMp3nuNVbfjPKsJOS4ATGAX64Z0Wwc96doqy0bXFvcdu7vfesB
tGWMpjVA1rA8XdiF+e/jaDyP7N3+xEqEfmyUd7s0HUNNG3chhv5akw3TSzQgCvBpbwnDGClXW2BC
haubyJ1a5iVBp7lNB51j/ED0enQyfYRCiWu/O4iWFKLDCH+R2/lvN9rFBEyScN3oh6ZQRCUAohGZ
1Z7R2nVHGSZWjsGPe2feIbR8o3gjhvLKwt8lcYcqcnLpcS78+RhlcZ2BajZ7NeuuRvvvsDM8iI2N
9ieIs3jOwJ+I4hHiut5rCiB1EGYJgmhyKJV7hyi8GwoZc+Huv5u3+Uiq8Aqr/dLw6jZXPTZYZ7IA
CAK75CoCVLg4TwRfEZTr9De3eYsFwapTsnQyu6LkDYPS+elMbDk17LPwCWiMsc5cG6PadMrsVP5Y
IwoivSNmpmtOXfVFzbYnnXtdrvSRCN1Shsv/JCaj/+BJKT65E362wCd26fKppBwVANm/mO7H1P4d
dD4E7rwdxPpDcc5UCO+IsR5pv0XulGdqh6rGVvM3tUu5RrEK//DUWH32fxEAp06o0ygJcWiKrY0Q
fUoKmMAv2SUQ4uIfz0D/bt9jcImtxvHPXdwtyk6Jp6tmkNJmp4lDo2XaK7QOgwu81BhmqsoC4Ozl
EmV4bTnTvVoKmz7HEZqKMi+JzyLWk4oE11XOGkPBMJ1uBQzHrXHAMMB6UGIOoWx0fVPBXW7wHfNS
MBnm4/tHeXyVCnj+lg8KmwJdLCIk5azdRuKeC+RUXReF/mujm6UMbx/t9cqPzhQxwtvgRBluSpOU
U7LJ38AU/aIWrUEgdZR5gRI2DiMUSLx2H/MoMnhQFMdU1NPLU5WDOyVz1uCnejMfAYfqiHvipjVI
EJ+A7XLTxbwSOoP2fVZMC5mThBP3Noq6uvySUDjL0QTPRq8m9Rwfn+lDOb5G3X7dHU72jGibTb2X
Tu2Ia9QZdVSDUuCfkEOplGj+ccJ3QcGmp1hhJR8mIhMygXV8sZ1qzWW8hvqj0XTxRHGKHnD6zxhZ
7nr5A7VI+ol2lQxYzJNkzstb8VxckwGxZ6BwZ8yr/nkTplLMPzkRgOvOtNnSKsYpSh5+g+A9fmZq
O0y/A18j0GZZdbtWyMHU884qYXl6RY6QX2IiLiMRwKKIqFHxdvEpP2KVmzyEkWO1v6pZXhzjrr9F
6HYeo50KfHrFMPBifPJli6saoHfxZgw5ZUS7k2k+kPqS6fPY0V9UjwCNnQVfKW6ZjKHuSWVFl6YR
bywmNOUb7D0EAOZ77ZLdO8XvljeotH7oFChK6Iz9i7u1RHZM3q7lUMHxNOX6RfPK3G6qDVpq00Xx
nZgM9RHRNdhkzyxDcjoGn8fwYXV/3Sat61KvwqXz5R1p36Pv5KTjiVvokcNul3P2TQ5//YLhtISW
zn0zGcMz8sHoPqdhjd6w6hb3ZMUuGt4mTfTJGsG1V7fBbmU6c5QEXEdfWzNKTV0XkfeD5Ua0x67L
zPihxfUSalMb48Mg9CtHuY4w7vFsuQc13dtXvjddtdqZAUwaTZSZ1cXw7/UEHMIYopbKLn0URhg/
Gebit0z1r1UoyMN1bbjcr2PhR3fkSG5HnMhrp4rVlETEChdRIqQatZuXNJxrfhcRDOTmYecGI8uz
M7MEvEM8SvX5Ph5/7Nk/GBSZfuaFcHTellNgdhDYctJ43t8LZdCSmt9aXJMtU9O81o6xT5FPY6+1
Mea9cAvEP6IE8kizQBfEMKkvNnlrYRYf0r6RTSnGvj6dWT/zrNrI6CbAWcSchyyTlbT113XcVxIX
AQqfyFAm5f8DCGlPz40eu7wbjbsJHq1jbXH5ETjxlqsic/UWPzuaIhs2gAm4Isr1OgB5K55WbmAy
aUK4QUyWStLrR33e4kUkz+wJJDiDqESST2CabmRTU3wAgOBtx+X9SFTnuaMpL3yWPehkc6CXv6Yh
QNCBsgEk4ySJd9l3nRajFLCiTFQR1SIr/T/XQJFemxihDYg579fftJjWEkDEDQQm1TdRs+/jpl0A
6v2uTD2ZqGGpsObxqszDCisZM4v3n5NTThUZMW73JAlYG3hBSkR9KD7Bhu2E73qaHlI4etqE1dot
BTGPIMlcDH2HOOJcsUwXp7oFDXqeoqMgBddfF14Gd5S84za5fClt+3ZqYj2Pn81c0a5emZKCTJe0
4uQ/1Q3+JNIQn2kAzjEhiuLWiZK7a4ZI8UWu61B4aHIcK1CG5apB8Gs4p+3UMQYdX+TdvfPfBx8d
Xts+GFx1XGm8EbjFJdYPObhnc3Gb9rthbk+/7/EnNsyYQpJNgaVrltYOfrcMmyNd0Od22LFM79Ls
oVOCNMokZ5vQ87dYm9Zs9AyV5MGinbrHiOu2wnwotRpa/p6S8PTmVfCbxSarly4BttBG0IXkF6nF
LUNjLtjVWLmNmJMoNviI6R4aD3Dr2JJDS4Jm6OJm536jYVSTwYN3sslkThuuOH7DfwfeIIMh7YfG
ntpeDxom3bailnWA6VuMxL49LAcDIQUVvdv63lXpO4tim8DoLO55MVqsl3ghOrE8Hd31p07NgRV4
Zi5lu4TRlV1m4j53HeL18vuAW7ziuslC7/rRQaO+Lt8jxHUWMo6IlTgp5ObeP+j/ezK/coZrhwOM
quxI6CqLKHGqZq/C4ngqFFOzdFbNLrHzS9XAOQkdvnSQVRXlKLEXtYMoMJcZr+V8s8a6AMLxwaY4
ofBdWGfCVr7GiuDV4dLOcTPtAWpxQG2/ygI5G0d81l/KnzEt53/OT0yQD3gX2UkzCEGArbH/L3pQ
WK/zwD+X+1LsXk+HOn84KWPifZYulLOmUp+grAY8DL/6MBv6jiR5W2AhkeTViUkgpNhdwhluT/V2
URR6p5WMK6fyJySIchTQ6ECrY+maeBWE/SwAsbNVzCT0p8E0LHbfGwubekkiwjd1xHaLu/9DU++k
/yD+ZuIcrrSwJCXTUSPXOSUAoxRMOb3z6sA42r0VMjLBNCKUbVpnD5yxkDCk0DspNugVrh5I9G1r
N0VVqlknn36m7EU+tLH1kshb+bDHKyeiuR68PayPeaXeV6WOyz4lUO/hByLXPCmiN9EvBTNJk2mG
bYT9RvDVGm1crrxMNGRCTvQH5KZ7YtOD6k3hqVSKPDDLiBElJzsNKX81sm0+wyfqOs+ML9nm1efM
/hlTwfNgNQVeLvcuH8aCk3Ji/tdFR9o5PWDS1puPvW9nYDri9+vBB/OzK0LSbdCUrGct1MV6zu37
/XvBqsh87Lx4y5aEDhnjlUmwJn4BklFy7k3RHDHoYfQ5iJXtWojbgb01kKv/9nP3AivekmBY57Sn
pgVUhT8isJ36gLQ+1lvA2oH9Q0VCs9MaiBhPWYhc/FE6F8sA7yzySsiS9Dg+6RELrkyfwKJr6d3n
nCPZcTNtilBi2duH+UrMI0jXENz2CGMUxCBsryOo+RBGzIE6puYVItN3NnD+dvkJYgjIrMY99h5S
jTmvCC1Flfphq9luhlKRWJWCk9GHrwbG2WxR8uvuyHNEkgQ3CzlkOrYiFj4jIqVq1nhPtoXPTnik
IqvEeJApYDZHnvgq6p8kxRWptUV1u3aSTYwWUfjDPt1ZbPcoYrDHdAS6kvzHPKMFO0Qsyg8I/JA6
iKxRxX4BPwOQR/sSEws4JACN7vdt7ApF9yBBi3PWghtrZFqokAgx5ycaO+00p5xP7cFBR/Ufyah2
ejPiYz77RDIEw7SPpwf/rdCMOkkVpKV7Ce4Mxmi6NnALgkyF7wV5m3Xi8X85ouH4eOm32XgilfCx
x/GEXdtIDdJhn7um5o17km1SdXGuUXsihFk27ON2Hwf/bbAfnikGf5XulCgl0Zb6PNOQYJc3jUpc
h3REQBY2hnHpxdO2B5xqnw31H3wBO0CVPEY0tcHQhRf4mRdJr9Y4LMeZ9xhnO4GRXg51VY9aNrzY
g91Dvbfn7mZ/Jr5zhugzuj089WNBMU9ocFwm+4h9X2deI8cgF7JCJDdbOQFMZADeJz/7gZe38g2t
Zxf9CLebD++cdwTnY3x1uXW0Qw0UqEWuv2AoL7gnN6YTsIHGHVdKBUvRHEXKFl/UV9f6k7Az/iXP
oIqCJBU+zJt+d8QUVzQgliksggVbzM5Ulwf8RaH6rgOrQie5cVMtN/UVc21/zwjnCVZwSfoF5FUg
6EyHJpH28iELc2Fz1alSIA1b5oZPjjr1b8BQqtWRPClQfmnYuhnVjYB2B5uTVSqt8JpG5qmdpdzW
duQfHiIp1lKfNsfV8ROfe6sFgp2wP5Fhh3iptVvWIKTOzjTSUOlHWNklyyZuur20d0HqFKozYwLu
ZLJJMmv6BlqCvLX+VHMpOx3R5yblu9esrsw+Gep7kqg5JzTVPGA2cRYSBUqIdhziqfxdurDtdCwW
2L2kNifJ2Nt06pd3GWNDRWREHFepxTfXRkn/x2sAeDNiqEmlX+VvkHq9p2i+28NMX9Pwl0UBCjF/
zzAIDsNUMoj72DVo7sf3FNjjaHhyC4e7nm5rVXEvSThWrml4z/pkKIjh/fkP4iDA774ialysfOZm
8WaxILn8NYPXiK8lcOllDpIM2fI6njj5Fx/T/qV0DXGg/QHTrgjw5ltmQPmVjSuV/DeTHD3llHl+
wFB65WdZYJ4zK8giOGfr12/Li/V2PDAhpBt6maG4EEr30EXekX8ThwfFdFG1JqPQBULX0d/Km4cm
EhvdRNFrXmqITGpWAMY/E5slZuFmRQHu/iY27sY18KNkdXDt0LA/hTKFMC6EXsDlgt/P2z5IE2Kq
XqxqQiSzB7/qmVwHXyMcq0dT2BqOvRM7+CIsOzBUdaS2Srlup0C7JcGX+ru1JLbiJyrH0OfP4qRP
sFAn4EU5eAcZtBdqgTCQoR4Y3GWdkLZKzEvRQTisV5yeHFz1RK2NaVo0sU/KUEPgJHlKx1cAtrhA
+oGQ8Tu0v4vwq0BRT7TrWHY6Pq/+YBs6INN3I6N6VxfJrvjNYG0f1vJTxG++WFZHSG1+9fwyj+Am
J9Esx+Hp2dDVkAkFEKCV54PN38kkW23lxLC6L/soyIoX5H0wq9fmcnYbcMOc5esqeAuRuXl0xiNq
+ELF8v9iVApzwCc9RCSP2vEUDNDN25bHZJkXJoVNWvrXc3Y7odPBlYEzRbo79B/dqgz03d3dGiTH
DB/dZe17iAHKqS1CnAk8e+ZSrLGdlzWJgjmhpzIcMEXfyyo8IWJoiCHyJ4CZ+hRCHzqYgw/yz184
Jpo0ulHB6oDErDw5bILGhHgg9jyHoT9Ca5HoHv0pHdX2HfIZ4dQYB07/Ey6QYX7KCLWvjfFEt15i
m81qKoALjNtRKtSa5s5hI3sym7inAERrF7rjWcRxQb+ZrCz46H2vE4CnYg8EuPBUaZm+Z3YiP8/X
Od0h8V/+AW7ocwK8VSDUXQ5OxFOw1kIGDp0FqQFzIyCKXJbSOn1dGPTJZQID1N2bEs+zLExq8yq2
Yx/Q5yq6uINGvCpa6l0qcx/fEirR9r4vmp9I339qu/oHefkqpTsInoViffxOt3yR0slBhYS0S5K7
urCjGiWiSjcORPyGbw1kXEy9jNTQZHKIFf0PBcug+PjKxO/HvgnJEN/jy6vW/XQQLYqB1tb9f/9J
LkLXjPYXCAoICftfcWTJQbimAL0/hxiMiLZeIjUTYMqkHyH5Xrhw0zjvsoZvdXbXdb7yXUL5bLps
NOKip3BKuF3Jm5mPvjZgrCpqLUw82oWTQC51t6qzF1x0u+Pv11z+daPBnX6k+cQhwnsKO8EqofUN
FbxpTc0cbwGMrETfz4RM8ehFYRbukgnFjkvySsugMmxZEjymPfQT5fDLs0hoqfmHyFbf9DvPT8p1
FizyBDToV/Y7zG4tmFg8TJCi6EVy9E3C8PdeKq6FLjyzLldidMBNIm9oO6npnDihFUxeZcNdbOy2
YeMAVrcbNGjvWalMFfQUGBMvU79nuyJ0+lp0eCLeY8LOj7Nc5hVr/mMCdsLZxgJG0MAJmhQpSlQH
Iyut201bB7pXUtbLu4dv5LwB0y3EixdiieunZD/asPNrD8/d72TN/0HIbAFE/Zw4SKKMAl5tFli4
IkSseVIJiK5668XBADtp+IF33ejW0XOqdAiaTWmO0m0pIrrBuNIeacDiuj3Sk0m+F04UTnCukCxg
Op4TmAndO7a4HP1wKdSxXY1A9cv2Cfh5WDnaToA8Im2hJGr87XOjQdYazF3eA5hH2EF4BduXGfIf
F8Zm8LaTPTTaz3mgIPDoPRhlLlS8c8mc1z1CkgaQF5V/zRrS4EDP26Oo83OPLjIdIE9jnHAGoJ3o
cO3w8s0Gwj+DNSnASf4A2yuGi+eDm2oEmTRA+1AkuGSO5xbUx7v7zAxhp4YDYmoDv6vDCG1f7/2X
aHzmHEuDyw9Nl8q5LIUhAf7/3PinHz6yZcNfw4OY+m9n/SZZ30fYDZK//og79HJbLuxLdxdZI6pB
/KKf3wfjkDZfeqUO+5YbBtLPHStgs74tC2Zx1gBz48SqMYznnpvuQGq1rhNdZJBGwybi8oaVcJgL
Fvk7FxLjcf9f3Y0zy9AeExOcqi0o4AQSkDLvclceT63vemE/Xmx1H2rmZb/2fJ7vvDMhLwau7Pql
FbyUHQaRNGAugibJ0OkhNI18iNU/rqukCvzXtrtTCzn+Rozx4JDYBzwZAc/Dzz7BpUzuCc+T8hOj
LDpPPE7T4dBdLPCsvatTj4yJaZ3pll8fomrKF7+7R0YomVsIqB+//k5MjAVJ9PjMSAKUmsFLgfX2
yWXMMioMbGzTPSMDPjqxXm/FhBiTrfl/hYvcrcTAyjQE+fryruMnuhiTw4LPGIvY0wCtShT3Osd7
qASW5rnvF7APi2jjGa4yE8mG7ui+NBdQFUi4WQstb+NJ0qZZ+Sa8s4g+dsqafiZKDCLWI2oBR/Mo
wlvfUttEP41q6UiijSdTKJhS4mJbvDMjQWp/7zUOoAZjpAeVd6/z8aGWHSprFC9oRJf6FkXp4rKa
lrxyLoByHSUav+/Te8L1KI0Ovm0SeR7XdxBZBlJKkC2uSgtvJe3g84wpa9NvlLktL5nUBp4FOcye
BzgM6hHnMKXPahFfEj3qEhyfQak3G3CoRo2v5WOs1M1Hh83p9OkrLJUSkh/yTcZY+iC+3RU3cbuv
/UMGkRgqT9JWFB0lIwAfDpaZqw6pX+Id5SXkQeohkmuVqv3odLuE7Oi9DyN5U0vZn1nAJASQtRs9
sgYRjXBlHPICOOr+EPWe6UhIQTkvz//jk/qOu1NwADZlDv+iXhwdfCjOpTUO54Zl4jcMhUtrA9hK
pg1PT31g/s/N7WFGuZRF5mhwHVHJ075BuLBhibMfB2Mxjk2QmB9UoPitiorHnJInhDlMQb8Gugj0
XemTYalNKG05Wwrqz3qEByxtf/FOEouCO3CsUqEMkc9nNNDwl6FvRv6QWudULm696m3sbEkMd4zn
pvZf7s4DLF8vXRzGHsDJkLnUbdnDbhZUQkmcbFs1HHeobjNAcK+K++Umsmzp0PG6PTm9FMNURorg
dCwCWH346qE8wYbq72e9s2K96gYYChEEkihHpFl8shleLff8pK53YWPC7ebLzpB+FR/eK82AT8eZ
ym6N38PNv4NtDjkYSDONGsrC6uPNQ25opUaBx1XW/Y7lO6S7GKYG2Xu0VK4QLCN8bKmqOpDJG3Lk
VR5FeWAOBh11BCHLADhXPLc1ShOkuTKJTM+sC4bCKE1r1GuqyrTSJUV3fQgo8z6SwwViTBxhCEvq
furyo7p4VZE4Xu+5g0QpkfyAw1Y3mwgudcjhVBsYdzLlRgH12mUwXiSNaUdx14lJlS9hUChwcBLK
oyV/lpjtMalbJGm3g6fbs/nrCI+aR4Wj0PkFYhrRVG3OJVPqF/8qFS7FVoNDgGHL5SDFse12K+dr
focfM/UQnMhUiGtz4xcDT//6uDnoeVZuOcB2fVYzVl0YP88bpx76RI4rsgYHowHQDASF2675OZ9G
zI7FdZOupcYF9A2eH8ZOYX1AdQ5NuMcZmpG6dcKXi1SL0D8QMVAlafYBMGllNmSIiG3Is/j6RdcR
/yhvPzrHnoN8cRiwLjcG9RmKEYT4DbbZSj7vvcArzTKwfKBBlwdjQl7C0/qxVLWCjCdzwfCI8ojh
6x5ziyUeIbbLn6CawGghIjLA2RgYLgyNqx0ULVw2gwjRP8uYqygH1sqqzsyP1eREK0HR9lJkd18z
hxunk7aCQmIqESvTXpynHFBryDv3ed4okUUTrVHWf4Zi9XVIYty+2VFGRP9huEQfPtIXl4IPf9FU
+AULvOkqK8iNVD0f4eHBVEkW9W0GUTQ3mGcnpWmus5KX47LjL3xePHtmtcaG0UFbxVGUM5zCDLIR
+FLAu83x8hgXDOpW1Oe8IZq4bPToAtzsqAvE2ZYBhd+pMhDIr9STP70nkNY7GZGAVmf9sy0v9qyu
RR58Zru/2ukTbY115H21KPOzQpJTmoU+2c7KdCmteXXRtAmAdsFRnXeRQPoj0KcDBRbn4ZBUErEy
H0w2REf7PXqAgLU/wXV98FGj2xE8r4S815S17l0uK1QAM9Vnaa/uwuB3qkSis33P936AH49rIDc+
Yofi+cbUX4/+BbkCFBUmyonlhQaN2kLv+6+unteNIi0v7ePo6hQTHtYgg6BgZCgbKA/UTn7Ae8Mu
d9rfx+iNTaKRHLP7QRH/jevSnX67wKHfpLz46vxJZb9FhX/6BnTdQhHh8n/ytzIsKnjnTGEQpIqz
HeVSsJVIoCt4fQQo4eKHQQCHcDqQdjG/0B9NLn8auvbBPfCEdKTp67BtHueeCNnmzzERLyu4kFay
54Kg6HZHob8qwHPdXfMFZqZnqMf+uHPXmpJ/BzNPkam+JIfYyUYL/dr4gRLoqOXWt8eul6DsLSNS
YbJLKF9g67+81JfuTh/TCDokHHUa0+qrAy31yhYmfqEsSbpdPpxf9GWFMhKkbuzK7THEOVCfGZdJ
pEyIynbXpJE5bJNo8d3l77xXTmQ/aO7H4tLtmKKz4wSaMSPGcQJDgVmoX6NFr9yH9TWuJp/PinYj
AohJTSVnYzxgCc6VcopSh5Y7qYPoqRZWR6DX6GoHSzDjPyp/wjIPAn9mkwHoRXwHwIts8rFH3oNi
b7Md6lV/I5oENnqYQFFAk1LcJMM4Hq1awZ6NusTwHhn2m32DcTE3punjgEVF1hjZyNI415x+Qtb4
h3fx+biGmPwHi6OHratQ024DKkA8ZLFeu3RktQ4/K+dWOyPwhAJunM3/Qk+0BNAhjk9ksGSLHAuj
NIWE5i7aPld4FNUR0EezXUMWFFnVewmStuugbK3NmuJgjS6RrIeMTOMO9Sk2Vi6zBqVRWwdotrj7
irzH5NeY8hgOHpAPHpkAQHwwfbqrIhkYd6TOS5BQFjiQ4CSwY92vbBD2WtgCIgVMfFmllR0jt+va
Ao671IBdO5LKMOXMVaBOf1v2GwT1YMwZ+zcTQiwwtE38JTkVnPdAYz6Zpa1Mqu49QKpgglOTlJDp
RzfwyitZamDh9f9bl/kYUUBQr/FJKDqvuRv84MSF9amKfnFw3ixlGXTZ7i4+6Y6WVV7bcvbrS817
ow56ieNysv3EoFXtO70BMKAjy0SFf2sJJxFGUBZqdyUimnJ/39zbcjQ/YiWvhvA+qeJNVNua0k7X
n/l0aajPos2qYSXO6Y7GQJeMif/JqY8VpLlKpKWu6L5Vckl5FkoByNeCA7EOZbV5YyDNOayInPKF
TIr3hGhvZFUczJaRCcRa9dS9+6ZOxF9OsmVyHEu4rvqrMKI2XUpiMkXA32eOOoKfiBPXvY09st1/
xL9N0bHHBlxJ7OSqqisftglClQyPHnhldsqchOgD5VARpqSyH4mpZpKuk6vdk8ox+z/OeKnp3GxY
nhy3XQpotbhweAXiKXfjHOY7+jCk4e1fQ76T+lIAFMoC3ZDTB8qhRI3did8nXT7XC3Ij+OzmIQSS
A/aO9BwJQjV9hwlgHVbdA/ZMsTGTBWAXFHnu4bUHgy65B6cpAJuG4ORwSsW0INZ6eu357edNVggT
hZz1821qZHrX+WgQhTTUSUowd/xv4kjUnLE/5KOfWGlQ9sNlDcnHnpywxrpwbwQ8DnLTG3wMW4lQ
g1xa7nVjVrGtK4M2QSb6IBBh+lwnKEwvn6Cn//NzwSuO7kajRo7kA6oIfumLrzpr7PrR+WiMScpD
XPdQOCD+HaEwsHQ+qscT/fh1/pT2ZwFvis+8qu3DSrEnqCf9f6tqlwgMiHqFJZYpnNoWgutGCsn5
9Q31I4wmx3oCaXe/vP871Okr1ul23t+/oHg5+Nw+DGe1zChbjoPU0sXSOjBdZMglo4/XNd9DcU72
TQG0RV1kS0M/lbI9c3h6MG5PqAHCrwv7jfJa+mua+7VATElTQgX4AUUhPkNfiH7MP2SGEJj1yTmd
ti6KmGsV6OSmVbPoNP7rnz/xOIl5wUnoIenUMp7Xy4Dzwbxj/U8wwJDbQVvfXjdbIONZA638MZ9L
FL0DGUzRvtgTYXCwZRTN8EQBez/z9jKwSONllH1MT1kbAW/F3muWgWY9r3jvh3/Z3rK+kK7RM89R
fmh4YJBphPqfBV3DCBrzBla9gaZ4npf+g+CSiGmCT5PopzqrkCPyLiFxcBquO7uALIPPLObXl3/g
G8QPLUA2pBpMSZXL4/pvSryKCZY96WGnASPd/MQLUGELLPijFuL2IqeycGKhSb4l+GYsJDU54WoV
pwk0INHejIsg4Zut4NpWN/xWKCIvRLehZSus+8HDs+wGRT9nOitkhwEufdAgGYk/ntWUi1xPW6Ni
UuzsS6nUZSYGwz5re4/UBB5qRNomodTKiuwNzTSVejaWpAL9oVN3BAGM72guDNa2Sbsr5W4EAOd6
gLTM5q8aEPJGRjjHcloTQ/rwi02zX8ZQq9/ls+q6OjytDKkZVcwXbDkWEt4UtMpPQ61x2GGyhE+Q
/H7c4SAnL4keDeVrkK1B0CGcnwIZXSlu7wEyllnxABe9MWDFdgWIhOtp/k+XXRpWeuoEdcoekXue
WQK5JF6unezqWG0ee4WXFUA0nGBhCoqmdZ5u3ygoieWECgAmGS516776/9rzRTFWV02UBvKNTC2E
Dbj0sQO45Mh/ZCmVRFUJ4YA/eEpCkw2+0eGlSUkGUWERyZBQ6/lsMR8d8AjCOIESNSZcKDI9CTVY
UOe3DT8XXVcc3SfNDw4dGFd5YRJrsnUxBY9OMJmoIb6EwuI7hVfFlNLG2FgroQu58ZqkBxRZs2xV
4nNCDaYNGNVF1+3xnwQI5+hNE+ktAuk7zhlhV5TbIh6qzN0rFYuQMfLzf7fnnu2jqJ4m6jinr2GE
czVBUpL1YzJMu9NIRx2Kc8+MYV22wZdQe8bS4X+FGJcRBZx/RggRzikPSnPtoCrmtzefFnSIe2Ra
mJ3VcDBcNLj4iBB59m8MtKthJGRxR8dX2O1fXlLdZFB1FnOdEQ2sRUTKII/HhFENLMZFCaNX0ZRk
Usy6HeBZK43RlBEaQASkUyDJT/gsnUrL3na6ZzXG454XBgijG18+gfKgGrfJ9q5CUGdXHEBYQ/+z
Jg42AdvmtWnvDIrviuw5SuwnvgqOytk5SxLRnCLGxyYwZq0F6KljTAR29LhSIeYv2YSwAxFCR/0j
Q9S/NQS0uwQwtA5Mws3+gN1njxqL756DA4FVcUikeeJlxYiK5XxiSLAdCsrmEws3ce7WMuQRXc7G
UxW9GQDWNw9K/HOFQzcdgf1l+tTJUpo7Xzl8X4MOYobKepZrMjDBQWBJ3Ar/4n7OJZMPWR3R7vwW
vbwPi/bSUPcIP/5eJfiK88rTudyEhiVTwXfNnsjLu5/CddlmE2daeOvOTIdAuLwhDrSIPFQ29qL5
j68j0SzMWTUoSUSrNySTtLlz+HODw8z6+HEgz23FEfQo5JoEiKgh1n1/qb0jM/iV95Qye8gWwj/D
7B9JJ7sIyd+N2UuG+dPBTXrOZMF5dY+g5j7mDhRRiqPLAz2Ilitq6zTJFpHK7eDKivmRACgNq3aL
lHizif3ljCXUKkHj+0Vn4u6H4Is8qQVRtiiR1/vaxQCQHJ/X/RFQb9z59h/zk3vkOrTXLLUpB19O
FjSG3mXAz/MHWiqWRh3fC3M+9jrWTtq6gC6xvL3zy561pz3y44FWUDveajZgYEXYL8Rjh0RBD63o
P5UYZvhSzdMWMrqpFybovwRLbiiG1c9QCfH/kcT9ra3glAFyd9ZXqLZQFNZ04sySAMO+x88Yhn5L
dz3C0lHmuydUDTTEPyPsjhkyMn+OXagHq5Rr5U412OUmFAvc3dXywPRXliBTAI2jkpvjNRV2eNpV
S25pMwFilPH+Ny6vItRAUDUYkhzqCxzZ0yrc8s/NduOTY3y1j8k6VtRzZX5u5LA6AqFjZgyhyJis
iBXGCLZ5yQKM5wUkFpcAyqZg0rbxAV1R3rRPjEPHyf0Yquhvkf8BFNikGTEIDfgkg8hBdVRR48lG
6b34+HHShxBNc/ww53dXmr5BsH9cG8LlENbaDFS5cTLuVMz8ZOtP7P1iah/j0XVuGHvmnArdKP0y
iPLRbXAB89bVVplXwd98uKXnhNZ0xRC0xcOBepnfJ75qdoOpw6UdwUVzif7TWMpDPlL0sMOZkwke
3aHBD1UpwARcaOv9raGmIDrNPFw3HZV+RBEirVMgfL05Pz8VPlzCKnJWXcXtukXUCyJoTboXg69w
SpePSZ9UEa6sw3WLv57iCuc0pixoD/LbsW1j7XOPNtWFzBSdo7kdgerzx6Ndw3riRPGHUU/lMMxk
HPfJsy8JtNRToqCINi9xT2bo82yrgpK9Rdb3NPfXOg3eX+aTa/7c4fs47XTi3ZhzIbcHyQpYDE+t
bhiz3jWp0hsBmt+TcavoeIhYLpMgYtdaMYEeY1mCOzs4gdjtugM4ii1WhWQw95igK1V1ttPpwE8K
nq5VQDflTVlFnMa54ScyvitHTE1DfXTb+p4n4CGP0k9hADTmeEL8eUhKbued6u4q+uAPYLMTF4hk
pyiCCdkVw3fNBLjbtwlvVuNX5eiGt1IaNotNe1oy8qAF/2cP46zJ7DAFd5hXE1+IMVOvkUYzLqJs
gFav2q/sbDsNFDmRXJD7l/+fTL8E+77MZqDNGHD2LxmNBQuuTlbY2kGp6orUJ27iIvKGK1tRhSWN
uth5rh8nBc9ViMMClcS73gV1ZT07kf70RVCNOsfCvyGHg99oS4K6gTNau2Ff/sQ7M/Fc182HBHGN
FJvwuAEa/6Rc3DixkvxQwYAsYo8o/6uFq8IL/ZVqBAwglAmyHPX9NP62k6OTU8cWZqxJR44wIcr+
oobRwU5m3yz0XASSjSgEtB9bQr+ynrp/d8ecH1ySwT5QovQwRh3pFZCrfI3FxPsRiOFh/Rlk3V0N
ijherSW4bCqklgstDp79X1JTJvQL/QUx1Cxp8qGmfYplVM7DALKl/wjl3ANu/tA1jz+jdlB1jkm9
ttnwb/Keg1R8i6C6sW/N2PGHwuZtANG9JAlzmSu7aOy0abYIC/DRyIIBqrEjLXjTkobfjZUnxIxE
zrTjHIC7GjZT68U2kDvRlPfv9tAaH2OsYlmzvDHauNDTefrvot1k//OY1aZakfxXfrY1Npzq1wT3
98c1iQlDso8jT5zi+px12y3taD7bAcOK93hGgcsLG4MgrDDOHkdSs1KF6NVr5xjmD7/k5d8eRZ9I
9FC/1otTlR4HrQUEgsQsDuuBNglLuKLpPTgbzNSEVfOfSha7fEJ5IK1cOeYG17Q7pSqA3l0racio
Q8dagvdzxpbPuyBWFo38LQSV2+eQ2T7idgJ8dx2FA1nL+Jy7g3aIZXwnMfSk3ktgi7L2CpoReFox
yv+qdzsKbdJljuSl9oY49fCqDFP4JJpQI3Nfv6Y8pffk9L9zcK1SgsUNA7Jmzx7j0fuNjiBO29W6
LFDuZCt/0qMxbO3z5+ao0b4Lqx2B9GnYhPPyz8PvIqd7F7h6BUSFuH97tzhbV82Kz8kSQcgtgogE
444kzmesEPd+zonJ/MRY33cbs4fZFXt83AlW0en8BfCJcCJfVRSW2sFB2bF+nehRIt9k8u0V52me
x8GSPyAmsPvt4uZQBti4s0kdISuffb7f6f68HxTGCNDsQcUCsbeJ5tdVhcK+iE93L5xgY/q6Nc2r
PDDvi3F0AMmD59lQCoaXM/89s7o9GMdD59LYqt7EBl762ijuJXkmn9AukQwCTzxdSU5cstm4TeN3
ZLx5hsVtT1DoLhxK87whXetd3AU5pvEyWgDrZxYzIBFkOOWr83g1Rmmh7PDONDWHCxv6mKOZv1f9
mmK8M6MoNhczLkCCDbeqoF78JhgdoOz8kszcCXRf3x/m32JhZJWpCdetg37t+GapATS+MiZAXh/S
Ly/yh0o+OESVsYtyvlKrn2D56gkNT1urNYqiqSc6NlJJ56CcbN9cuB6LRk2Q3HVRFm5XRHMttjnd
zsv3nO/jp//l0aVG4yZhZC/iiUjhD/blpqt9KEosLuvJyH1Fdjo8Sn9IQHxZ/7lPw+IahqgP+wIt
0pvI13LXuH9sKwqZGnWEpNqmGRjhfV0rKfXugEAuwQtqHr3KIwJQ7IoyNH2ZQhlpbQgGH1Eryiya
4vZDiPVyxDtuaBP+bvSABP+tK2O3oKW1lebrJGARLmVr/s2TjUsoSKuJauSDSa33cSTY/b0GWOHX
JbDeuUb42IWq9T8neTbHODgXpnXbOZxCrRJMv5ScZwj54zxFpnhy3CLdudPqiu/cIlfOtBHdvYnq
y30JafGTXpQ6cQcl/D/lg8VUvI2T7jAl736QWSIILLsMTPTgOawtfQgCFZGPWoP3yH3Th3oNs/Ym
wIjsaWf9vikZ3RWAlB19XIIjnnUHrU89YorHYW1EzIM1hqaD1mUhVSugiwtquP78FSqJd7dRSe49
QTjOqP5H3MbL1CDgxq11ByeBlwy+qyzT657lwAhUAIPesS4/3UQI6JFI5kVQtvc/lQuXJF10Xrls
r/6cbJ++Q55l4VCePlDOt6E/jWFyku0reo0icN5Kq8k8WOjk9vEs3s1o4SttUdxTeXf1UuATbevA
r454+D09i2JfRyliumQIK9RGBFbfLl5r/lEXYXOOJRCUlKRvETDqoXAjsItKZttDhME0SjX1WgtJ
TX+nCl5GDtF2BajH1lse83PXi9R8iMYRlVSgzM2Z7QrXY/Ygi0fww7EDMrRnoPOAQwG/QBCXFZhX
BSSW6X3a4X/URNhymPxqtpZQjOirNdZPSLi3pzJUyl83ijj0TTvmlzsWZaBfa0sSC2y9LJUHMBpc
+E4Z/96GbSrNpWkBFg5jnddssmM1eKJpK7vQkLTkNwgBB/7DRDXfhhjQXn9eMS3ruXS3R9SDSYfb
ivYZpqxZXjAHCe1quJygJ3vYH9/D3mdsOkesluKdClcHnnxY5/YYPkomdOxAlSZ8+6UsISFosww3
xxVOLwfRZp0GsqdeqbyhFiF6MruNccKGb8QSEzk8GS8x4fLjj2u7/27ZbN6bp7hsSpwwdSUtcKk4
FVDFRBU70lGefz5c7H5a/ICYoVZOfr6gop703Nf7JLp4fGArnWg4GLcYwBWmcvDIkLno/DHqLliZ
7ulbpntCgaCAYN51px2RMf8r3f3E3o2dNRELnZP33YxDoeCoJ3i+FYHxcF8/V1PUnv0ApslGbf3F
4fdTPy5aQ4ipdbwYKTaddVTH5VDYLIC6hapkL7RAALWq8DBlQGQsabZd5dLlDFLmRQKThUVpelmI
JbM8kzoUL6QpLP6gibRJZuIjcXrKEt3D0q+bXGj/p2tAiuuF1mm2OXFoHIbjBp+OnJaVbtO7Hs5M
ab23SP7ZWUZQ9wMwP4dS6l1m4byIkN4ts28ViG58dvcVQltReEdO8v5ifqi1bRXnCTgrs1hApDk6
VcHs3Jt3dwHOg69DNin0tlMR1Z1QAxvYv/uDOxq0sY3MqijcHDGjNGjv5XT3hu4KOVbbg3AyZri7
YfASuFONjZ77j8OGYzhwXwH1h16EK87bC3u+XBTpCsgETh/G0vae6GgBChCPa9LO9Ix1l3NDdgRj
eof5jb31DbWEU/7wofTdQQ5OXPEkLmcfEzPpUTZBjANtufInpPXNg4QXRSxMFiYf7hKtZv9r1r2s
8kVWAHb5FlRo7ma+UL5j9riPAcoNtrFglYrW22qkkEecfijaelTqVGSuMAfFctwzo3W2GB4yE1E8
bN8N/QZsDWJehrgY/WoyJCfg+sB1q5hRVSxfislaJ+VHh/9PD35k/1uvLXhPbf1NYu+eWdpqcejd
wAgVGxZqqTRXf0dJO5EfXc7WcZlbSWBVSk7JCILsHhLz3mqArUfECtUCfw0lov9TcLCMgqXPUbYt
Tj7ErSEJtsh6dcujnIFgT99RDvY/ShMZc6lEgoDwyP4zDAwOYslxLeiYniRXHhZZZa2LyOS4lcuT
dZtoAVF5r1uuI1375qEWZw6l4jBgsV5eHKPD8j161QMase/yh1ZTChvzJTBO8F6go20XLehNn+Ra
BAhcg0FurdN7li7+iZEXaNKxGF4GTsLPMhLMtkME9WeRfVxAJz3Dga8t/YffRIxh2XgVSFZwDxRS
y4Sq0GZtJFK4qrQ59g/uHtkiXD0nD/Wx5dYjawgS+5478Y4Q5sV9ExYrCmf8YtKBDY/JQClNakv2
kV+W7LZ3AZUeO9TI9SkIrXZUjKZna2yIyNPFcIeenzGJcnfTqlwhaNoxzHDzZe16b3LW3X89yeY9
Y4/YhpCIOeTnUaiuFWrGRBxSeWvo2YzjsBG0aVe3ZXIeCCXNVD8REtjpt99u6VSsrHUmXhk2Bqsd
mP7Hl/UrJ8/u3+XRFOQ7K22MfoHay6PdzDyTtrC7PVUZbiOcvRlLgwwNkj0TjiXFfF5ej3rrhgug
gXA9QHEFxKTsybUWJE8vSyYgGrOt6LflQJFFDLFQNq9HzcfLa6FslsvdlCFAplmFzm/e0y6fdMm+
Fiw8T9LWBbWWZYEhmmg6alo3C3aHylTSX7X3S7E91JhaENEbukTwTCb6p0KzP24+mKC1VvgM/DNc
NhWx3nYJYTWc15+D4xfyW2T0atUun3oivoB/iUCBgKVpCzT6/nNCTWnZz2PPGmhuAE78OhMZEj4q
PDebUfq9nivbTUG7finHQ56Z6a+q0DFM2iY5IMqTrSqayzgF5ST+bCsqNXbsC0aw7bEPx1WjNqp2
1LYGz7Zb7zCeXumOUACMqAblyv/58VNiRqywxZ6e4b93wZZ34YQm8SUizH3oYeh67lHai5LemBmx
4Thtu3tlNK9hGq90Bm+NhLCVFl31nrfmzy/k1nSm9ExHbYVimBoB5W8pWONLeYUDQmui5gcPIP4b
Pk5yCzV4/7I5MnBcNxDKnSOoiU+mVOs/RJqYEDRH1X69dN5PpzdJWqw5xSSJ4fB6nYN3HhspFBTl
FiXty8PKpkZLP9gDFYlJSnOAgDtJNlxYrA3cBAprXOU/qe8q/7c5DKFA9HSFoZO2GR7gsZnJw12O
lihNKMIOQiGvJuHoBDZnfz0296ZLvEY0nNQjo50c42pI9hitMJ4AVPQX3YiZ8Fa+FbMhHyvJuoRQ
ntSWTe2sczsSQ4e6J1qnzQyHAH3vcBGhTcPnQOVk+fW1Gm8prLth1zqbcXxZ67kDmb/oBpnKL8mb
tBsYTgmdFz2cJVY+qLfP9yoXB4f6NN0pP5+mWTuxZzuXltOmuUHIT3+uk1zWRaj1OzIy84RokNFu
AGPp1CZ07XNN4E0/1ZDUtEHgk7n7MpbmWhheInkPu26SnxlKvGuPZeB6bWleDW1wQ6QwbcUcjhne
2R9GRkO5YHvUVcDfmIZec7hFAqJY6JUrePoIwcox7q6IMyD4BueiM2V9yoKRyiRSFuyoMBMHRR0c
Re8f8W0qEfNHC2YTdgIZLzBSeuJojVX7z1Qk0pXG/uzBwTH4mbwd0jrwLeWTwZJJJVVXfWe6DWxH
JNlvr1C7td2cEk1meZ8Nrf0hvfEvNy4TtMbw5jgELEU22jyBo1jwhWcilBQ6o6kdo8enJHhUg7VZ
FQMaV/8yTghYkcDnoF2oPx/yQSlz4tu6KK6dsCArWjiioZrXYWykogqtNEdVj7WnSOeBemTC10YV
jaWlExn6GIP2wYPTfFgQ6Da1A8iX2rfeIeiTv2JBF5neH/3J3uJVTX/WtcOllecVsrsL5hWtf9MM
sBudHLKcHD6IN4WkvO8TD/5DY3QTxjopiGYbeexQcJdiZNrFKCay+SEXZLfdsVmckYmj/dprnjrn
LYgaw1FSQ298KMhMtPZbGHUrJsuJDrgGqgsldjTFmGlCgHK609ckv/c0Wd+NzJ0iSmFS6HS4/9M7
u1QwHB9sol+hHCmlIPeDK6bNHKeOrwzHEOXjKSZcn/hzSkXE+vC8YjAbH/Kf51SvMsXFtBl/ocvx
/mgYc8HoH0Kgrj0xiqnKyKnA2wj197anoyAHnZaCmHPNvj9h2Pzpo6j87Fytmx4ou+mOBdijGfxv
bZyYm/kvn7MLyOAoSFXJM8fZsblV/Pspo2JO6dvMXjmzIoP77Q5sCgh9GJ/HZ+Ax4XpTejmGSHiN
B0NA6Bvs3M4n7HEFI2y/IgRQIEyjc8KNtRD/zkyQhZ7gJ4ZD4qUfCVKUT9Bv95co4ExbYGnP03xP
C12ck2rN6ZQq6IbLgbHk+D+MZqrKYEssSinvobSBbXLG5seQgDtME4zOl6LZdiW4etdjKM+095yf
E/OsegdpD7yx6d5O0mheO2QjsKSrQukn0hBczC1IUt9CmkzRBuCK1348yyAVxHoTyly+GjF67rIz
x1Td2Hqij8YhDPmPqkGsF2+zi8KNcl6Ahs4q6RHW4vbb2shITqCuHdKn2Q1kfP8V34Xd5TH0iCOM
85FKyGPahQzYh2XD+AdoklLj/K+6A/lHzwIsh3LRGsiBkWQV98BPlppK3WEdIPYfrLFLE3ktapNA
qCXAdEr/GVcdAop9fd88LzbWPyu5bbasyI64tS93skd62oMotrCKS4WDPoZf2xBYKPh7euPPnFTL
4lMY/HTfp0eH09PAFwG9UYDpBNrZ3BNydthuB1Bm7b/1dNucWl2XArTwnUtkrWJlAOtgUmFMMnXI
/cU7m018FZjjnnvKAgDgjSH+Cen8jJV2YlziQu7PahGOaI9EBdUe2L2LKjh5tAKsWMJP+yiflA1I
5GGdeqrdFfVGT1cFwZfffru+Og0DaIV3HjqwpdYzGySyugFZJxVai0ehVH/hcpP/J+2alCUl84Ox
FTXiPlZ2Up4Ku1zsIbWUAp89M2kOlBKavD6x8bW9QgTf1GQW6oDvtOqYiFLkJWJd1jHg/oxNRckI
s/XJj3nqVdwnX/D+yw+HTzNVtFl0QxSmNfQ2KkVRvByFOKnWyeTV2gKmdI+uMijbAaZga9/bS7m9
bKDUAaNdPGO9dzilKINgeHBi0t26zrRWl8ytyYvuqR6WQ+b4Mt8t/mEeHTv8b+SRuChdBaZ/Gipy
tEfeVgKIhGqvm3GfMCqwT8/i31zkYfqLYPC/eYXKV4odDnaLAz5Zi0TAlz/+xljY4TsQ6dmd6d3u
aSDU/LGqM3aFmwK8qerFb8nITtJ2oIXIya7p3qgYD233WQYZz+AAt6kgGHEbWTkcmx72cq1ErRT1
1s7qzO6SH2mzzmQ6i4GDEb643aaIFJabl0D7MkX64O7V6hF/IbmvaYGGfhGWqVpZwuxVG7wKbiWZ
jikSscrRK+ORELtF8UfAsyhjGjMXen4U4pqMxJ0yW/Uhy9jxl7DrwXcvuCKKmlOmF5q6xC/+t7Bu
HR/qHvFiuOY9z20N7/au8lNYQj/dC06zyB59iPsLLODpwq0O3A3QMhFg5nY0uaktvzz+JN7Xq4FK
jN8vewE5rzOXOOrYVY110mkqkdfG78Bgt7CA/O5+D41QzOfDtmkZ9k80QpX1r1IY7q/KA5t4PlfC
qgOLwEHl9NQvpE3+IwPV4dvYveeYkqPaI9AwoJ+GUZa56DO+rXJVet1hB9mGbRucDs2iH8SMBMg0
FuGPhJosFJS5z5pIhJA8/kDjbHPiA8c2oiqvG9J2Ss4nPHVjOc9dqFIUAKPFqO32OAlNs014isRb
pE3vrHAibxnaDNQLPe37P9XpPgbFLmr00InwwKMtckVAjabot/suOHjpq8unbc9RryOL7Fp/TOHp
vSuR5gb0Tt6JCKBy1JYf5Sx+XQoODDqPkbtkiTZ0YPc4SZPVD5g0U0bZemm1yGkNltMAnGvBF0Sd
Xb/K3S9jWZ94QlbKjZkBa03SqH1SNeV+2/n+voo/sEaiUlHGJJQK/K8EslPy0mVTli3YOfOn9HxU
gKf3fJorPdx2oOxYRQ0Y0B1vVUJt/yGkf6VSnMhUfbP0CZhxyXDysMy5lp7XOzuLhgp5k3VY2a8K
zsX0rDcrI87y+V8ptEmbfCf2qWZeX7zY27p7fKtrIBVCBt5O/6M+A/fZR9e80Zlt2U9C8HZkqcwU
GuA7TzPKWqze463kOIjn7qV1ZNBV3CEEHQ67+NhEVT3J3cSmzp/sTy74+fmOwbz7GobL/Rt0QGyh
gEAYaeTjpeAqyyJ51VlXMn6vDn2Ula14ynfYAkyfIz/2jAx0o7Spe1l+zei0/T2Ld+HKmfxAMjTS
JrH7M6dPvm0bCWEqiCdqxdRwJdGWFn1GCZdYnlKjjp4gMsW4VAVVobxRU75cOsaaiq3VQ6LscW8q
WN2Q0HchBNUY202f1tpZlzrJWO8woCRVFyXTqITv3iHLRzZLdOht8Xdl/vVSuZUtyh3u1SIji78+
04udkD6YEH+fVVB5CbEBYyn1rgWlkg5iBioVWnzFd+zWZXVEH/x3Seky2kRatR+Xtae7ZiMUDYJ9
1nM+7TzqE5wvG3ZBdjwK8tMpd21qR2lLbOct7Ld5JvvrJ4hx/DwHHQkUF2N9aDYGpBPJAHX+BT4V
8RpoQ5MFxaKyImOg6KenPcppvUVpl7I4mmxGABxFV/10xTcySTVQDb5T7oBn0/Exj6kTogXngp6F
z9a6Z6IJlmNXm2YtwQEnyyyO5nPqyKvEU59vlUySOq7r/AQYzTUy9ui1PhstCKI0HqFHewll4jRV
Z2Ac843+RP5YH7xCZ9QGtXx+XlwVEWqk+xQ2pYJY9q6V4gHI0etW5ZynCm/T6fNl1bdJdovzs8QY
Jcfl6Ty/KlgZVG2y6z8T2oGZxVfeRjdZrnR3+jrKTKF2YxIhxJq1V/gK2G/WpZwy1faScgB85MMj
wTk4pa2IoRWetTwQmIfJ5rDzMLw5wLJQzGRbvGeD9qKWg2x6W46ygKUTqMciR9KZ8shrGaiHPmKY
3iy/tOS1uKGGbjNF8vBrJ+JQ3VEHvXmGq1H21edDzeYFHcnFigrzVvRtyMLXQSTz62z6bO1uAbKj
QwRyTNwWdE7CulPqjfyUofvNvwgJzrDSVLYiyPyeswWrHcSnZ+ogTAOMTqDyRc6e5NKJGIGC/2hg
GQ+5EEqHbY3FGzzfKja8gMQChKhKV698iqjuvUaG3Z3ZgpcizyFqv1U0dbWasOqM7V/EGLyYUK4l
jKQdb0WW3lQDp59T0PsaPO0OZkS43aM47DM2wTv6JXnUdWxgRlWDM49b+BOf0BAx+/0X6r9riwXe
g+sEDLp9hTAkFUcOMY07KSBlbYbnllqa03M1Yo3LFu+XMyVdt8Y/vyktduI1PnyFOJ/jxZfzgGru
4nwGLQJGh4l60qD8w28Zut+UwvuYtqStYXkO+E8RPEe8o1Po29WTq4hSLS+cI5nj5+SSESUVe3xp
3u+nWLmPLsp9tcgR/bx9bPSFUxzB4Ntg+VGThIWiuCx1RpPU3AXR9iOKxmwHJ4pal84lZQhavehL
yUT7cBbM+bh8R+TW9xYwYDvVa6xeFxKGB/0+pOWH8q2aKdvlkbwaiDkoO3Ng21rkUnDn8ylIIQ59
6XBzZfsuxXowYI9EECtv7AusRK8bJ/KJ8/jcTSFji63o0JjsdHdHFOdJ/e81QCD2HNrohk16GOfC
6jqKxRbyvCubCzFj+4Yx68HPGyzgAasHmTxMpXgPZIN2sdTRLtQMKdoV3L6QZ5Vvk2OsUdSx18os
qQdHn/+tISIhlVhUW7sFwSoJtPMOMmiCgeLXw0ot1/89QED+E7Z1CxG5KnYIZRVe3PauBS9UG2Pj
3my6de76N8PDTiimTh78jXQKJBLTfV5NxWlIVdmgd48hUgNC4D5UZ2Ed/W8yLDHow/Utkjgjs8mL
PW9HtWjmWZLSBWhJmidEPAXzqjp6ULmt/H7nHPG0Nz/lsclOuVER4gtG3P4AEMSM1Ba5yt2sKQqx
ves82lxqrrRKfaO60r5yXxgmlJ9UcSBR/mqB9T6gi6UyDzfhLQwD4Lt2+j0rla5orZp77+rmoyKc
zJxcrpDfk9SpA8l8smrvCHfcH5LY6lSy0qjYUQDHuwEvquEQzt0TD8FjjWPdq5l6Nvm1dgzn1GfS
isycHXriwum1lmCm8pKIqKdwDXrgBLVHI1EmzvmFUp17GYwZSC2fn5v0UcdIqMCVaUTFWheSZ9uC
f9BdClSS+aJibnUARSlidzzjkEqBsSnsY96VgHvFyA1v60BjNpaFLehksHRKMnunpW1VJ4M5Uh9v
m8hWLnHoSdjU14vIFNJDuIvOdRiFGbZB2z3WgGGFR0mMZuavMi91DYvbUCKsNtv0JktqtErECCBW
NTVrTfhK2PmiEwyM1Aa0+foqWLB01lYavCV6+eQ2l65TIzFRaY+a7YV2luUzGbe7vlwWWnpGRabV
e+hR3tF/GZERpJVHx0W11wYkdvnoGO6ZFAoXMhZTRLXLvSAThZDn/4XeEhxThGL6/YwRZEacnQnn
ldKJSvRvfMiE4mnxdCvJ9KiwRZZXaA3Qn6Jhgr0rQkJhr8XXlg3Ak/d2IdrO9mdRUtFjIdK9OntP
LgcZpPJg7csOxB+XmACk7RlM+eBYY+HfjexKkXLNOVxnnSOjIExhk/a5IFRgeYn3A/xZkQ6EzX7s
oRRxn8OWLTdBDk3xtOub3D5tFPiShbTkK7UQSuo79sWaZ2hANw24F2t0re5lPMWHMnHmlCZ96Y7T
/Zqc3mJbYrGrdjMRSeoQwPSf6/kPTGEvrhXIuLUjlvPPcb9jmaf1KtGiuaSs0KJhHHPB+Zip86Y/
mFvU0q3ReOujK6iyDqgv2g7jz+ljmI1ktRFgSs0Gwz3VAWTGkgzRZrktFky+DZE+gCBjOPBQpVqC
e7rVKUB44sOF/fQtgJK2Y2oDmQgxALVttU/oVMWxqemCjpB9r558+o6eX8u4/kxYK6V+A0LzRTWv
yI8ZUnpPKrS3rzU9KgyK1OqaCWIntiFil6ty9TikvanDRGLyHVZuzvJy7Esy1mC/+EpFI5mPvgy1
i3/9z27Y+Y534+PVFovcIRfPQNRXS8unJuXRqm4jKkM+Fo5RrGC8FPrFDXvQQcMUAqW8h6QwVNo2
9UU9GwWzBjSldlCw3ymrRhMh9EHuF+OkeX6gQjWd84JGNxyoa+6n5kxC38rQlug9WnjWLQKSR5fc
Wf67C6204y3nCv50JNVeUQIMKpUd2H5dI6j+LQ4DePYXjmqOoCh9X+SgB9A0Gjg/wTRmiOZK0v2x
uch5UsGqw4yQ8JhTQhyx7aF3/QNpCOj/VOgAfITBFbqehajsbQX/ZehFmkMwgeNlCneL1ES8tLjg
LaRFy2XL0JpXU/WBHD2ni7Uecp299JBrTRQ8E5AXMEzQls9FF0UX9wxcTjJQEy879R86qS5T7BTO
z3f6U8xiXTwdeEsmV3lZF/Cqpr79aIf57SGPQurFAWCLY0KwZZ4JzYBG3078evVb4tTRuKKjS1Q8
2brGMttybNFfAw5rEG/W9fk8YFmIxHHQfmysBo3Q4Xv6IRvIX7uG3LShS+DqLpnyVHuOABmM0Q0T
eu2Vqav9EY4u5LdRkPEJ4rTuG+7jv102xNZDGXZFXsZ1MWeS+aSRPywhPpfJq1MwFfv7yJ2ahQCg
hsmM9RxD5AxbJI9z5TNPA5D7y4cGWo68z6nlMzO6tWXLgM+HZwIZAX0PbTBxL76pUdI3HY63JKFB
DctkBkECQZjbh+QRaLeNa4/4vfWodiKmGzwyIp2qjJ/FU7xDTMZXYisKHb03IzXbZYgFNwB3Xg32
oBk3syhT/YN03qmiMTA62AB++Yrr6/DXbwtC7Yi4WE66E9/tcMNNA1ppfej0alCWGB6D3Ap9lPgp
RBBDdLnYC9bL2zML9hPNqw+m9esI03CcGW1gML4WZ1ZZl/Xx6lBx0NfMLEAUjrswxSh4i+giWBU1
tvcTsKgREy7OoxULmPn5G4LyHOsZqwgWtQhc/b3BIAMSm2oh+PLvmqhY4tqRifWmeMIBmgA+VMvv
bjd7cl8Yckfv+VYhY8DQnwK09qQC97hu4sk1Q4mCnJkvG4VaxIuyq0v+ltWIANYpsisS4MCUt8UW
fGLd/3x37DKAxIw/+qvGUxT48qr4hOHPDa91qIfsRCS7o1EXhVKr+FWJ8qsOZuFmMRoiV4FBcpqO
WESxNlARuLUXofD97N4/G5u7XLg68wCvfrMJsSgH/vf65ajgKNTyzqFZbCblXpVccL6SJgB/dEoL
63zjj+wpFKYY/NfQXrvnkJXgAbimkk9/X1QGqXw+wCUtjg+hGNKOUIcyXoniAUA+g5RPkq1z3Q46
BjLh3OS89fkyLJ5J9x25hlBB/mAGKs4ZPLZ1RGecX0POQ/ZdwjJHpmJHBSrCEHljQp/VJpSZGuu/
TGw6GNHEUr5/YVl5UUL/KjnXjhlPw2AH4nIfGXYTUis3yQUIQnaT0bKukw7lNXDfmcvfLDBK+dLl
O0YG4Oi7/4MuQrYlMywONg2q2fdR2CrwqAy9orlORn846JGy7XuMS0BYABBdxqJ0z2WJ6pruVyfl
PpCTeURNbmh5X///2xwFLajh2dmzkpq4VCIBy0yMB480GCTt/IX/ntvVbFzarRJyCp9pSP4hDCgt
98rcOxF2+rs+7YrO9G8fFJ13B9jfoEgTcP18srJ27AAfTCw4H2xcfku9dcF0iaSSe6m6uTFmV2AB
5y6b2kxhtXo3+x3cpLD0pG0INopfKbcciDmLOtwncv8d8be7YBrZpNimu5y6LWQnkxhZtWaLUxae
9Zl0yjb/jc83/PPa5X1dYBajpz8wTN0iMaNG7Mptkiyoi2qkBYuIGEf2DckgE8C/cfCj1jipAkuE
Ti304oZGq82/Y/F1f3dUreqrUTqPgHnMrQEh2CVvEHG+CLBgDvPlRRLt7Rws83p096m5NXKoVX8y
9DbAZytm7Ov7v/vKIoJn0FVHgcEBxOxX2dACv715Esx2TLkH8HFR7mKvlrdr+4iI3QOLDaMRYAMp
mBR4latawuCbXvjrgsmYTvgy4EltrFe8fNrH8LWFQRN+bkkqO4Fl3aL4x89uzYkScYAJR1izkKI3
AM08gbgww6ID18Kyvp6CfdixRsxX0owy29YFJgaFyaFORnYbMiGFsE71b6Bjy5GP3QwVs/bSFugF
y/JHI3UQQPJ1ssfN4hXoCpLV0RVpQACT4PPqp3O8+Tcv5Cc+Y/yzaX1kj07eb0lSy6J7DLW8OIup
FQK5a8tThXt9YTZUK49z+1iZcchiYGN2IsB4sRR4fSF7JOZV6hNFUoDQ875I/7cspid4dXLHrbX6
MN/zUmZr+10F4umYus+oFoUv8cw6lB19MDtXcd4EAN1AVkzZ23nEL6HLEqLApgrWlH4xXuVCzIB2
sPYWrZkW1lqgkbEYswfjQMAXWD7F7WlQZHYWrRYVh5/5GQIBy7e8geoPI219vwpHgIHpCitSgPt8
7bsnCwo+vjVjBsxYSR2oi5zMOgtvGU1IDaoyGy384o293PxS3ohxUufDUTR3vGjfLVIhlPVWvMSF
q8/x1MygwlhPFBr2LRYdJJjlbNFOOlXKo45ftB2tBQGBGppylFrOyVrfP35svPFWCOKQ4RbI1x9C
yho69xU5VhO3hSKv0nf7EJw+7GjdDHhO8HMbu7cdd3DcjDtCtKeMwJhlG5OJISS+GqytbtEOqgs/
sn9IS2I5iRUJGK6RLQxGDzG0bgUyDTtpN4N9PkhMqXvwVijrclabsI8G1afBs1wWNgZrmOmvhsWC
ufo2BpDiKuLZw23NuB4vDGBjIe3uuh1F+QxTmkFhRYhDmdXbRNJ5T/kH6n72no2alA58FPMaM+ZC
szIDXtq1n8LKgnApgFQerII3XE4hNlUb0RxWJtypsjqSPdA7A2yfZr4lX0rcEO2h/VJbMlQf3KDi
YaT0AYGfhDM9gSJS8SAJv2RG4uPvMcJO+Znx/hnKPolE60bm3eIAbifhFKxsnTzEbgwh8yJAgAGp
TXfMrBbeX+XN3ICnP+ZPBSQ95OEddxlX2kRW/7oNfGn//ftOuF0Nt3lN39/TtUveQIKbJ1eVCiv2
gyuiZK8P1mtA38SZgwa40d7LI0qElZ+u+4ya8AuStRJkR3dmmFLIBF44LSU2w3hW5pO0fdKKNVfx
jEyP3OcNL2dmAoNaUOqqZMVC8PSAekL+YJVaxuX2R0to1kp//RAUS4I8Q0vcmbXztQjhYiwSDJYZ
Zr5FQE9ZdtEjJMRiynPG0lpBOjgWJvFzCi6I8yTUZgL2Pe3CGA4pqvaXQxIBqS7Gq5eWI3LxZaUc
lxd+6JMWd4qDwAMeYLEwaoq3NqWvd1LTR6h5/EndO5wwlcFsvRFNvJu07sIKeyHKpryI+wi6c5KG
GtQX2CvPAD9pr2K9eVHuYEUGdIztcBR0iXWyl2+on9RDO8dck5syxDofPhFwQaAnMmkICDR59a09
C8PhNJSjYVaOjdDdVr1VUTdeEB4gZSwntbkdW8vFQA2DhUdxBMozlp+0hsK/CIvI9GrtfEIaOXRH
F6+Ef/fQ4zlIT71s7QUMOwbAF47RwJSwJ7Es/E5YR6rEoi9zl+DgxOEI8uNdZhA7ZZ7vTO4Jz713
/xvKwE7fkmRQhiUr7d2Q+LtSjav9F+9b8iEVq0mcWnqGkb1FIqA4TltIF8KczkGx4zUcVZj5p3lg
M/G8PKZwof3o2gLtorLA+WuTLX6bN47o/IRAWq5aQUrB20YDbGHg4suMqz+hRYR24iT/NrPQ+qNz
HDhg8/pzaDaamDyWhxZqDHAFlW7Z6Gp6Dd2MhFOlQYqXC5L7EKTftnvJgMtaSQSIbw1FIFDnSD5R
8QpyAANHykB6iCdgl5aylI2nuMAsDMxjq+dAJtXA4n8dyhI48DaF2/qJKuozWVv0BLEZ3DFcG4RT
hmUuR8Zgfa/Bulcy6WQAktrO+9rgoNci2CLXEAZKPtWohUc7FbKw0+FkKWjQq498dyCMGAnx58Zr
MpnJKMDpVXlJEwiHtJKhH7YRq/PQrfY6rvIBcnPDfyw+PNzt1N5Vy+/cZB/WCRl60WZMT4Aw5Vay
iesps/IaAmaf896MNWY1MtA+Dc/UqeY3N9qZAzoT+0D3MlnbAd23QKO6H0ouOjVm41i4tW71VMTT
Q/QHoxDx+2enDU7vGRwAzl7yXfaWoJi8ynuUQzx2owVcYtmqMOs3oakVo1bUc9nlBDUewo540v2q
ot3DZAeutoYs9xW/I2LskhW3q9kEPIo57N380kOy1Yiym9ro1mC3TmUF3dy372Otkrrqa8NwIp6p
TL278JP5b7jHzEzt2u1fT5U1IjxLXWfG5DHlCgjQ5VOaWNkQowQAwoEc+y9zDJHUXEuLsJapOWw5
ecVeL5PrMC99a+s1Y43fmDjGqHkL4SRSpR5ihpJzdN2Fmwq3P/ZSApagg9Iop0ITiNVNlF2L+cPw
HwJqZVDDIKA9k6KkTA73Mx4P2Ieb6tDS73I8rsY0a0G3xHJVz9NgwsHx2XiTHlLuRo+m0ZEr/iFe
TjDjd1MGGhmM7s8ZUerJmZAQyHwpdLXTBjSnNyMl0gw0Rg+kmqQL+UVh6nK1ErOq36UEaUN5h36I
B+1fUe/mCyxZowJOKYUbd049a7b/FrheYLfdGDns8Qpf00VNn5qY4FaN382D9HUtTqUdzyhOzbU4
XJ/5voxdtRQ7dozKaeJPRtLYwG2S1jhrYvRvd9ikB4GOYJAOADktem98tmJvOFmgXG996aRKFW2b
FmdCpQQLeACgMt3Aq4HBStyJ7UyGOmT58TIWUjYZ4pagMNEqUCLcXZJ3BMJmoykDMidX1g82lAK5
G6hRuFyzOQxrqSMkfzLdDyMbkYlJQJyS8jGPNI+y8j+Lg3hgADVutU6/G0svGebAzJa6BQFe4pCk
kLAmZRjT8lAlXzAlR77YC26gdLVnZP8LS5Y81dhalSLRu/00Zy9gNF3w2oJFLzFZRTmNzmilM/mg
m8svBuZ1ERVMzIk8IJueDG3BltzVF9l5c71eUMimiPOVyVaMju4MlNgHARrUJ/vHHPEvFZnqLOKl
zfMorkYoLOSXNaoTnyr5NYmm3It5sm8HmDwTWIwMsZr1MOaLe/uU5DPd+zEIk6cL0qDPUF0CpOli
reXl2NfwUncHwgt1oOywGTKOo95nQbMRt3wKZmwv8B+T4rHlKbDeCEymyxnbdSnZRp1a0Iii3mhQ
mv+RB9EtnN8yLy48OnpR3/cgw4P49nNsgpST4vcfRUbO4MO0mVDRCeB+jO8aZOLEdJ1dmEgD4H1/
dsnHfhsPgIsIGmlQtAnMEXxnD+y8JPgnP3mmMAFg8MExwWR0lb7xxZ/lebSCg3NMO9leLXkjt3+R
F/6Uof7d6c24KMSgBZ7NUg5HSAh5kbT4LGnLnrOXM8dD+pSpUR6e0228Haa05G7SW1wIofH5VYwu
NBsTTyi64rkaerCWjaxzybDNek9w2bygtnuUmANCS5o5H2jeFdAjO4LNgF1ZpE0IXZuSUXCpzuFq
5/8HueL5fm+lNwdpclPBrfyM+w2F1oP7O3DYpAnIn0TaauQxeYrMc9DTdEj8n0O7U/3zAi4SuhDT
tWvOw3SCz7tlLp1JEOg8YFm77+yyCJc4FEu5uttrbkscTgteSGwq+WZwcLLGyz3QNBXp9DhSwkQU
vzV4Cx0TMOc1KCTyljzK0+6FSphQv23Twb2jCDG70X8jB8XjRbVz7s3hv7kbdAl8jdw+T+K2n/VI
6byvIqUHiszidQdQRjxN3fm6w4U8bsL2lkpDIWqT2TxC8teBbrXs3ZhieV//e8fGbY4Lurf5YYE0
7UOE5tE/a7ODtnguRxWXSo3Bg2ZkbWZYJQISXjo42PhYNAFD+kUf/XezY+9MIpvQkCmdsIaaJUfA
6FRe7HEhrMIV8cFho7cs2kQLdkPq9FsNX8JpE/dsYcANcvEKvnEHCclpDUxU/lUVW9NUnp3P8qA9
YzSaetJi2sdMlgEADP0/CcPvt3WmCAR8eKm6Y2oPHOBp1KYAFp3WhSIaPK92mZ+0Uhw5wT6Y6oaP
IclYYVTIi1AHCwWm40jkRAg9olDUMWuBpUcgB+8U5d2fJCeyHDFlhk3yuEPO52FlnCZbhs0tjPHl
BytSif6z3d+38ntFp5YkvG5fpFPDjRT/7bzKeQaEym/96H795iwlOcGisSLGUlyFlUGadyFzItzs
WIIg0J8LhLeHwC/ZhQ5aYqgndngmPTXYpOwjZgSYYHJrnWzyS1FbsKu/tXBgJnv6uolQrApUmYvD
JaOT2FT8Vjs/sPSSuY6+pDRFlYyhAK9oSI7L8OmjDfWbBQ47GKlp3bblbhhf0lO37AsrWXCd2KqX
w/q9yvJJsfc47BQ38ff9kuKHD/j9icHJ4A2QDdGzaZgGlfCPukyLN+mmzxMssWsR9csmKhm4Ecxm
90AL8HF1Z5MnrpnG1/rfKbVLhTf4vJWJP8LZp3WBnVYeD2q718D6piEHrlFoADAMEKRnbUOR7ePZ
Fe6gfsUzUQ24uEMTMPsqaR2Zgf5L/TLV0KcepbPsjMimjuhP9HnyZEWyIQlJQh+8H8cI8rtZ8LhE
w0xZazILbtClEOYj9j+k/l9VY7A4BNxZhzmJiOKTA02Zl9/aKNbVCpkrKohaFPyKb5tQxkvBCZBp
mat+IjkEPjeKpUihQDjbpuOO8AFCjKRR6NGhfUGBfn6U6pL9U0sBPEb0BicQfE/AIHJX9yLZo10L
JIaCmunjuQ6z3T3H7yqfw1INGyb4C7GD0mmWlwz93QPyQH2pBZGG7C9rv5EpUMQpvSC7myOrQXgH
9k6BSTGqSjFY6iTZUviDZWEWCsFZcfY8uTEeewCbBfUl5IqO2vRrXLMb4qbjAsTcJTEaedAz3thT
zLUvHdKnt4UgBmoPQDTO0PCN3T3QtbSgjVz68CbghXicteoOKY7T7GHQxLbg7aAvr8meTRSYAFVW
Kz1M10HCKAE0zD71KCavRscrdEXsuFLvwBUtmhnkg/hbgbjvZDaPMVaFriRwB/pK81N8OPWvTWHc
DNbc+peQoD7WpADjP50IkOiKE988scSAwH/urwzril5hdmzjYY6gZ7D+Jw/Pm+h8EWqvUydXBXIt
wk13XD9pjD4/SyH9S16GBmVxHTLFkqC8v1gtfrloeQrwR69RVfGRXOdwr7E14/W8zOdRunf5mDHE
njW4aeATuR2RmVOBvnUJBzRg/+x7JZ4swYG6lJvjjtlbspHjwalU4Dr68iN46OIo3qID89KhWQvY
3Lh9XLzkH284LIczCutWIR4ojUV986tjl6MIpbLmkOY4xrRRE0J2kkWzZpsrqqb2U9rE4GMUUqnx
WxCKTZkMimZYoFlVqSaqtFr5WWAhJYvD25h0ncYzxJd/Ihdn+y2YvoRrOlWIqhNOZYhDkKBgAHSn
tBaZoypmMUar/c7Jzqc1Er805cSqTNtRMt3yK3oY/AuhsVr/T1PfzOv7VgXItYikmKx0+VfDkwq3
tIJkOdwygcWzKoCn7HcJ2Iw1YAwtskmBCCq6Pa35vQkuMbKdB2DQa1oCmmJwE0qttgdLtNJnJ81X
nl8gwSKF/bOfqBDpzNvpXfeg4+dmtTcXXCfhkDoWOGiK5ONQVo6F879dKdUtLHqhYK3H67YY8x2Y
qhIsC4kaPyRBG5TfT+RxneYeM7CkWp3Fr0sNS3s53UVHHlHrZYgneA0Y7d2vBogjvwxxcsGLU/uc
jjjhAue0ZrYfDieC5W1e1uKuuGG7WDB4G6J+stcuaJuyIg674ZWgqPhwgI0N01lKoHG9O4gtfbK7
HAOilRdLEYt+Q/tni0/3B6xwa3NK9Jn+mas8bzp4rE4BoWfynJJpSOrjph5W8iZw6rUHaDjAasIB
t+bVPEVZay2weXR6JblPjreMNOiwRz+Y5fL1fXrb5flayfr8ueWS/CtTj45gsxMO0zfqoiB5tcrs
i7u+W76AeAORLS8miEyMOa8Gm55lx9ijF2aQ1seDMQlZnGLiPZsZXPc1ksVlgzd+FopUAHFLHnVU
kBDC0qbbmNZbcm0Itpatr7UVDrW0KSBgYakgLkiTn6aAO57Txb1Lz9S2JGN7PBnH8a70n/EcdP5D
ek8qDkJDzKFlKun7Czm3/Vjt3v71Kmspr7IJyVrKMVmUhe37RPwxFe3b6EhzvGp819wjX/8oPla+
I3wa3jLyq5ZzaHEtTi0aMl4jzFl2c0xqvh1mTA2UTYTJlfrShJX22UJA6vGh7w98CFTpp6Gw5en+
QcMf0ziPCtdfmxmI9chfj36cccwnxHbnv9eEo9y648M9LUADGj0lIGjIj/J+M12TkXwV5ppecmzf
M7+JWbEbQ+sd2FDyJ0perGQIU+n1DccqvMcZioDZuA5laN3ZqgMF7BKWRSJsgV74fMzbMW2awdwP
rlzkU1NzZu49JmayKBO4OfFYAK0MaAJVmrJAbPHalZ7OmQY5R5W5ToepBA4u54ESEB6XQ2mpKwgB
1H90pkwdbRZ/Hiu8/SvNwb5W40SImu+QDyMBq9OhSdfiqFsIXQx5JPNu8TYLVFgtfb51wqma7mBD
2VXaW0jtNka0TGyVVppC1+0IPPUSL/vD10mf0v1UdLTAHRhyjqfWRMWj2JuzfDlKKzhnLXWbEIAm
PaeWrBcNp/InqG95wf0zdVvE1c4vuhHRbgxI02bSnAgnpYyeMgoo0amdDPoWtzlrtCIATzW515rW
b7UCObSZ7jWpLKVit9pTHoHv9uzNZIGIyTwMm3cfveh9FWkZsZW1FMaAFTVzdwSAGDJhydFUeV9A
lnoJIiJ3ZKSlyum3YLvvsO7nAJE+WGHYn/hLnPXhukEiN/DMbPyVLUbIUCyeOyIBlmfXcPy2gvbZ
mwv8MBWV5tHnAlpKLp5hCPpjM279RZjnnuEaUABVOREfjfKn2MI8CXZlKkWp7xTdtsX2m07W5HWG
TIK3A34nwqx9Rjnxf0lpTgPD1iqQpLuHX1LiuhyzOmi+IP8+6M0eVsguO4azy1TGqdYvwz+hmlc+
16b4eqTIy1/pvzfObCH0lDPlRsnvthYenoXP5lUQdCFi+az8WChDjIYdpGLmVm0tDlEezS62fy1p
otcIV/3XKmC2Pv9i/w0pUFQC7OOtWIj09v0mGg1KApfAvMTyXSFJVWKc7yKmD2vEtRkalJiFGEf1
n6hugBIsVhbkLIpGlMJLd2R67CULUoMfwiFAnJHZwex2wnsQaO2fHnWahDGvKga/Lpos3G5+Dyv7
54VwzCJulW/3p+B2rY2ZHbV/ge58DSsoyY8D0XWh3i/pz8pwW3P6iTyooWYQ4VPeHKXYZdHyH1hz
KI/O5NQZTKgKu7Yrv3YjGZ+1LHBzNxNoe9liBDvcJ4+3IPkoc5UWDgac71jyz/IdMNEUUWlnrtrJ
9chcAq7fpB/hatKyAPUhjOGrBy1D3baaWKLPdsf5atAocgDsrd4wZA7co1JA9Mm5OyfDq17nFYyG
FvpykBHujxfMbASAnVQvYK+NgjyFYNOEvgPjy2TaFCoMVR1U9phL4UN9BMfG8+Pu/YdavOAX5PaM
yBFqpfp/WzYbG/+MJsveXabJHRfHvj+wj74By3VJKHM7U7f+Gl7oBCaaImIUAVW7lBThtPVsLHPE
N0MTytk1ecogfugzIDvQlV0Ne3bYZHmd62tRPUzf7oYWxBwDqJddZPS9PBp4vsfVXnonOk4r2Izb
uyQ5mynA9xw350QJdm0DPjQXy1y20Kqcn5xJpjxTZ5ijvVKiiDgMwi2JvmA19gzUfq+jpEZEaR3C
aEk6QqsyNAz83FZrSfXGcbyltOaukRrfQvBY6Lvi5KxDul9y7lBNARL4xoDkDksRy5oA020yp6N7
Q4HTSjO4umR+l/1O8OuyEDpe+dBZ51oFjw/x1mO6y22YIDu12unpW0jsgm7vU9aMB0dJ/UMf/ib8
R1v2q6d7tTm6nxeUifzZRdZBSZYj0eiEu72Uze43xdHw9gfzqFXu+O7X9SJSljMzIMCMsdtm4HIl
ozqiPl3pg3toPdza0Xmnz8U1uZhJjIPM5sBqGeIhZ5sIrXRYGacblzxxoYGoI1rXgr/h9Coy6vCY
7mZV4rsOw3M+9kZWObK9x+eE3lWQJWvHe+rmY6E7yS3Wh2Btdr5QXhWn+abUZdynBuNS2ub9pMVB
FRwXKMa4XIAlkggMvMdrSzFJ4vcPzvYEyAzjuWZ/F25GZLtB1qsa6pvimA9vjI6aeE1aOgBOa1Cd
6eR1MgmMuWXKGvmHdjIhuFk0O29wHb+uldomzkvwhadPi0t6o4lqFgsENvUyHf+odjUa8xINUDvg
7rwKqhEXKTZHzzElCJGlrLjpRsmPE7uwu8NvXE/aQdnDkTh9vO33sxZOXgkUSnm+NbnFUHs5BIdg
QtF//beda8eP1qOMJPLgkcn4CoQNDl7/h0F03K6Wz+9Rjdyd0dpT94LwCB8vFTLkjoC+FpsvFnzV
ssope630m7/0HULiixewBgbgk+HY4fcvFaGMkYyVo34f8STLiC6zqAfp8diFOpWmCIH1RuMOd6En
3BeFC4pVGbTqxPmlsbD/OGNfkNuF3zCzaoF1TRnKNwIf4H4pTSLxjiv3o3L+XeY6FyfxT5T1sM2a
yNvBXwQ+mLNC70jsDz4rlWgc0USqbezWqy7S1iijr5I5OxkdZnaEWUIeCbO7B7j80OdwVhpGTvu8
UHwmdAqt50uDFqOMEBwgdzZbcsoV+z3OQLxlGfU9DXgMMAombEe2JdoPvDOTVFm60J7qwy/7MMHi
YneBpv/8IF8Aw4asfUW3bV2V6BFuYiahtPCJtqQmGLD3p0CwcOoLU38Tvv8/BjsN1RmJnD1EuZAc
y0zlSGWHVT7yQ34KJf0cIBRZ7MxP44G7O5c2jq3plCGT2fNbM5t4bUXPlzQuZC1EzWl6ydUX2HD4
c4jxtZZic9E5SBp6wTmzK3PuD+0a85BGKyfrB7WdEkCtJD7l8T0C6Pel8SoRsFdpc35vXFFqdKIx
3TQXMiRcut+OY3BKrJFaVxqWjsdJNBcx1wmSMaNE3kR0C0W2A9iiJ0qftGc7dFiRma2ynX0voEW2
tp9kT7HcTOjheyrQ8orjwxmK/WySn8J8dIlWgWwh1zkFc0CHlg1rgOFh0ytT9UOui0xW2BkoaTvN
rrBYkySs26VxAXPxIo08sg5XKSF+/GMPK1n6qO95qFB6BPKkEbKwWckEXQ3kFV7ic57q/sgLfzlf
G7wgnYKkToLfixmb/Q3HUiwpbrD9d3Hnga8q0MX4Wsn3lD9O7lToImo0Gt0ETQgNOVXMq8uurD0l
/2mE53s+QV+NdajF1OkUaX2YSFygg3XYEFg9vceUTerKpgbJIRrjUj3Bnc/w20eakAcGbcrxakQD
06LS2wpIVROLEtbxc0E6a1gveAgkIXOXu2j3/7v/bTD9wA2+kTkRrNjKZYDFO+JJK+Y5lCPxVBSG
EJqFWxDU27sk+DV0M/lGHFO6P08BYIIKgXRXdIAyvrVptrRcgReP9sqhoEbWRA72a8wyM6qOkDAJ
uf1ILUZX1nwph/JH0aQP0zcsC1jjw91dEc+AaBQWPXqcAcyGtXcOqL6BSQJe0vWYuQonEDRr/V2G
mvB9IHE1FHO9TzK7a4+h17vu75E10q474gosKR9ZrJAtAac49NYGTlC+EqKxPgg0CKALUHJ6PY5j
jNlNlskyMYTCMkDzwWHWzgiDP9VvUZmOFAE5SKyZuulE4iKN/+e+voN4A4nXT4QmhJMcyXJmymua
76FNcvE3XqoqNn0qPdvM3N4a3BTf9uwRYhK4FSaI9DFX2lsLHfWOHvVA8OFsJNubPPHJJMjoqG+k
vu0Rhrw9CsWVzAjDmk3lUrhw34Fg1slJJyXMgRSNv7BwtZ8QF4lka4dgSikm3cHETmedGtPd8tls
tY3nay00a+Mq4I62lbQAyWb1k5E0MV9e2oWx+6D9yVsSfmFwAoDF/m2laKztrBpMafjOZ0QhksoB
ZHR8NYX6DoTbd0n6c56/Q6LvqaCPLWSkVZs+5Sb9wGYdwqpxb7UkffaRo95dHBUMkoQfYLs1659r
psvEvOZo0sTYKo4U3DWkKkC5zg/u+SZvTKdTQvQ2zlR66eenu92s0oJcn+o+4dVd4E9VAOLtHpSG
v/7EqcWwdgt62MaXlmyrLti/UZPedEIs/JYtMUqLnevF0PT2Iz8qDUFZsSKdD91rlpUbP/gsObsU
WzFgER2xRpkNWMelnuoOW/VqdSrqDUw6xX96/kWjTPCT3pj3jPvSvmCoXXkUQXgrN2vAXYJ77N+1
014rT+jfhnO5PPbCqWOjhuAWzA7W/8dmWVlbv2UDDdKRsA8XWJzt5Em8ZB0HmsUCP4xPDCvObgIz
nr/snPbNKDD/tx4Lzj/rlYa+cEO3SFqI+raK5bx21OSnslUbwhGV2I+KhwD19eE5pylGAwJPoByF
AvWDt4OAzeHXm9BBjNNRslQI8CN2jQZ5s0wRVWApoQ1SsjSTNSp3ylT7/tTiT4YpSJNqikoOcT9N
qkRzTaKoI2ViaCVrbkh4TFKg76AOaKQiYtovZXO2kibir60cEWjuagDnYYoMxLBfhNx2nNevkVcG
U4FDjwxQXzDA7VHIo4MN5K2laRwMTPpCbT1rNPFWZBIkYnklbJP+khtFqCcFLqoDUXHeo8jCJkXE
DuLyQvOjNYCNMmjFoT8lZMIgvTDTibzFv3qW3su3MCfSVkvTArEsAG3e9wd6vnRTWKylNOdBVCKI
Z7ksUyNsaIIwjpKXjNsZzoIfHQzs9gtADCg4zQrgi4XbwCNeanYYLX/vbZIJlh1GeHuMcjAgk4lR
fG7RMndi54nQu7XO+bLLUOesIZVpNM2GqwSvMGZ5z+eBpFaQ2eYWvh+3FvR6OgVVVi9NwfhKcrFm
k7l/zDFftpIJMNLI5nZvCYbdCsXxhFC1C0JGfJvF7s9daxNy1HzLoubAcLAtYq/5GqGLvk/mjqVe
9Dq2URFEkBXWDquS5lzQEbhkjbrXPBX+tjYgmLwAUgrp2L9+NdAj03HTpO8O/tZe1BZSaMw47tV1
wxE074wz3j10i43EUiwSSTStiBowBXwR3LqqvgS2CqIjT70Dn7OuHc7N8qTlPyUZxlTsn7T0R/Qc
76bZbQh83ToWgxla7Jym3mbEPELJ0o2wBoPRVUHya93JGDxYgAv1tkRIvT2DSMpKJ5yAiROZLo64
nvAOC/nlDyZMAMEw8z1ZTflpZXMsE+buG+B6YS615rmIeJtRLvP9wA52Byfqfuf5sJQRqVX21oRX
ZEIf2q9og86YAqFNJ4Kt9BkENQp9gqukbmvBbPNz13ezH1DMLzgyhq2voUBZxemchYUfihNm9MNr
kn1AUD1H83dYtJ0+Fy8kkQMong4k47KA+/6GiqJZVaMRNg82jBjNFy70EL0T7GEagYnBDNuWu2i3
BPq0Glk7gvX4MsarcTJFDA0u+T9/e4gs2w8+hcfjnFEaarcQfX6/Tl9m21GB3RdtZeCBdBt1kW2N
oocMUHsxATxZ2//rRqe+40jTGr7YFOaskZdPKO9SlyOZ10f2aGbn/SXzrS3dzza9I6xNfYC5cLMD
N/pivYJQqFWIcpP2hZfCABVYCXjMXljVvYZa4TVU5F4ButIXBTHWXhnSkvZjvdt97IMkc2JoO8Wa
qzSrLWC6CesHG5gRsHAlswwCJTzvPkXU46Qy69BiR7IS7x8Bz55pF++7MxWFlBV1Ky0ISNDtpNC0
/0xwdvJm5VYz6BEQImUqebrQMCP4Y2kvSCbrYP+anfS8VRQBdnesaXNwe85ICn/ZVVTn+A0LHN2b
fKJ034gYpdda/VzHU2880kokLAdPhE/WGQPOMVfND7K4eFr/kpQ27Cq15YwV27hfs0Wqf8tsJWtS
vLae2fvU4B+YkDgzg706eR8x+OkhWeNofjqDJVXcl66RLrK0wsocJxu4fHoiF2cOBd0P7GOsD/wB
7F+FXiVxW69fj6qtOZNnHprYdpN8j3SuXNFN/xcs2wtxcVdhydcoI8uNbbdNl6Dz0H2Lq3Fm57nk
tdnuHoD1pTPzpFsvL0ZSZcD4PqUqHDw+pf8GxXj7mAHMJpfiFuXCg9hs2glwBe25n5bFxDCk4kEv
DmGGjrFOZeN40q8TjCOSdmvlSpPRqbWLBccVdgdaUWrq9Deden/pv+bezbXcxfH665+PNl+6+yHY
uxtlxR4OE/GZ/Rdcf7xWWwCcYUw+7jTyE6TL/xuikzRRPCqmiZC1KPv5CxuP4NfiL12G4Zuuqi9j
1/al4XpeR/bIbdlguE8r0G9SKnk66nkKmEqmBwhCYx1HCcDyryCo5eyhoehHvtgoij6mKeWKe6jz
G7wtKXgBPtwVWxOUo7DFhSUhIJgcZ4bx/yCSlMGk+4SIWpW2a8uMzeXBcBc0gARDr2TUX0rUMOZq
/2LciUMKBI2q5VUYtaAmJwaPXpwxzm2TaS62F/Dk9GsnC0D4j2jIRCQV1dcmAr6kcTNL/m0AKNdE
WBa8uzXgqYcZbBQb5JgCaz5bORsIig3TeMQcuHqJv2KgmmopUIg+L199vFqF0Wjj2s9Wy/sE4nhh
fM3LTzl9KP7oTarFn0hqw9y0Bz6ZtseRQAwl+hDymh0SfU4npFUTRetN7iEFE5VV2HCbVRuB5VEz
GORIIfj2dRNhFAo3LK461wHfGzBIcGFyDafKHnHgIqkhXXGKO5nOvx5WXypMpQ5rVCAlzDen2yBS
JYygNCMRIKvpQ8RuhGmDMnLrUG0BfxZU4VYJc3mRiO9EYaDl1aRXV8/MvV22u2jVnYP0/aKDyYWG
pvxie8ewMa1z+E71fCDu+CprYdbzfIn6/Jxs7PbvSuTGlxfkCUz0Suts3vudCaNbQZmTRTgbzn7n
l7Enfac30g3R2qZIBfVQjxPSl+Uaq8AwnOdHOok3F99JXiwQRKwIu4JOcrhOAcMQtF71zFoSoyif
ubZJ14kglnAq9Zk6wD5MSRUmgKLHtOq0b5+gDWfaIt3693Em+4Wtg6X7TdxOvsMykFlzeuGjxDPE
NFmhZuBjTVEkSxADLYwyAEs5cFBp53I/htmL3IPEQi0Nnn10jxEIEEc8My3rnXr3dWsFaaRTqAo1
j18OAq91c43ttO+IbDKo54fDaAAnG+9urKBYD34GSiBjDto/EoOtmaJUo61qxrG3xW7d1TnTjJY2
PIQmQC33/WoTlshXs84wVPstUKttIfujbuFnwXmDeeD08ME1ix67rsD7ZZUxc2+Ju/IXBek3AL5I
C4BuJekYB2LfqqluH0N34qqnc31fBc2wOEgrRtZ3lGLDWYEHC6ejo4usyOlm2eQp1ek2KSYPh/MV
VDNr40/rC4pWjygY6hrkOU+WuIafoZ3wJXOsxi39iMT4uTJ4YkIYnc/a8U+IUIcJmcfZJlfVIzc3
o5sbdztNAZMxZlJD6Tm0Ra0El4K5iKTpL5V4dYug9JlNS01zVttMPY25z6QjF7sF8fcHAQN9CmM0
Kz6WpTtUm6VtA4dLYZbL2MKppoG7WdaUPjzZeXfooNO9dJjpAoVLGU5UYeOBDrl2bARWVDEXK3tk
Zth0hQ1UY+h7Hhh/0rJIIJpMabelqY8JEXszLM+fkS7n0FmVd/KO6dVyJaT16U2jpE353h8xZvAk
zZWSW0OOVzs6qXEzFTA2tCgZiI8Hs0oA6/b3+roF2viNvB1xBvjVz+fEIWff/PbveKEBkDFgqveH
1Hy4HMldn03lAtGJ0LRKX6gwl4JfJACu7+xTT6mT/+vH5OGSM31j7lqiZFUOvObfrwsXIKcJHAFt
YCD42/pGmNXKXW9wAogXfVvz+X/5Hlcg122YVKhIRH9dfHUvDSmH5Xs0AvfL88PH9x/AHVI2HvgC
oyou/359zLcKldPjhgXfYevnHp8N4E1dpzcLzMBsQb648n/vMzXxWDQrQuvcsKUgCzxjK+ZVWBOh
oSzJge/dN3TQugptGpWh2KNk/gmKsdXFr56gNwJVJACrY/tgfpLCltmZj7HFkbTSRQCHRwQRssRC
x512jzzqbxW33JPCWrfGTZ7S5lfWP8dkwTyN2wv7U3FPvAbUD0UYUf/bB+BDra5/mel4hlqMXAxn
UcKtYQekHeEOPGsfOqawMFoYcuy9+rpz8z4ojWRUs9ce8ubGam10Y+qk5RFd4zO95XN5sviEjUHL
Urz8xJXRD7wXWB+JxZOphdszfCEpi4cQxQbd9Cf17VwQSTgF8rSKUF8UPsVbCqgvcN4dt+SxNpTG
ovjQsQ8BrHY1oLnQHrfpp4pJvCX12iNAtBMexr7ZtWEDYoAKbOTkII4bZOfTa3VeJ1alpSkzovwT
TGDxxce3y82zXUSnggj3mRM2iqUwu6OcyH8GCg9ZfRJcn/+qAJd5E33dcBygCGFiVaJYcJ4axoHY
+ASd3jLXbZWaIBtWjzH9NN8m7bJsE0PVu0FFElwh760ZxKb5Lpsg4vUT0pMk7jjyatXnP/qS0/iF
OBraBAOLxRlm/VxdufInDyDgoVkHY+rhKJGqzzpa/kNm64fDs+rCKD5zKlzSKqJp5mxC+NE6eqjt
k7mDShOe1XB9kL4gZKrSMwPYg94jpedElK+PY/idaullU4SqqEgBsYFfgiYgdiPZEpeNIqf3wxED
pubrcE/KSWVlGWCU9wQrdBn/Rdnz7MnYshg1JPwcfxSmnbGhcbXW+ukQdfdec7jt9XLF6493IPN7
fTG4NqzK2BxjexBrFA3X1VF6ShasTpaTX9ifyX99U+QWnRm16YS84IQPUmpolUbbSw+ph80ol9QH
FQ/u1M6jZjo7cXMXdhe+OzNBH4Y+wBT4cTTLCwdnhsNxZhXk+hqetGzKSZ234blzyB2I7yxaXbUY
kKxz2clEwDK+cJv2RcIiHam6rC2m6nazer3cDDbv6zYNzZjd4rbMJY8VEroSqjr6KfUTBEX4BCsu
OH/fVuDTdGUPzQrq7PUqL1ufX4pp7ZHTRwNRkYF5frF/7p1mVjAzqCen+Dsu/d3HxJcTxwjPkdZo
SWq9qs+xMKvLgsdqRgnIKAId6KaCvEYue7lj3tTn67uSYaPTso9AFkkbNm4/v78ohJ4cjxRRuTzk
RhP8C/lqb5IQaYRKQfbzz1yVQER7LAbq+JdabknHw3XmRTOVxVtCgKSn4mBkr++ID9ghVfnhz6z9
Mo1+AxY7qdluphmUi7cgk4DBdC0fthfirGESYugq1g0sLGVf8opfghq4ntgKIsO/2hgODg6XgqQw
M4Q7peu8PVpGf2c5wJgspDZMRESCqbKuPjQXG3kSaoNGIRjDfBJiJ/EBgNm7S80f57FJO5pcjLyN
6fmTGcRZgrMLpRLy6XEwT+iPrtZbIsHGhUvnQ7JOuyr/gPphCXj8XuzzfWAm4GgHcOIvUXeCERjv
aBlB9ZoN/1Q5rgj0GZxXY3pvpO7G2lFKBGCgSsn1LUELEoXJDeKytGMvAE8xmqVMsY4Q967B3HDG
V/dJ51vxyK7Pejhs7zGtcV/YBIIPUcim5m1KronTJcfcu4ApGRMnQGyCI9sI/HyKGL8Va8prqZLH
j5Y7GQpfTw5T5eM5CNTWtlNEoqlK8aJfHeGCgsmgevxyTldAv/wVhyRM8/JcSnLcYDX9sdYna9n5
6XRueRhw0e+8IUXinRo4ndQV9ExGPjetXJupcfxvfWVpIeJhdkxazQ41nYFakpoBffl4IuNIm69T
hh1FWPF1ZdO1NoICiGe5GuMKpXhZxnlbe4QC56wWyTybY75mecRTzuMELZN/3zTv5OyjLaGx7tKh
NIPbly2m7nZn+fOfpoJy5ALoJ4zFeAGuk9gLMeBeV75fVI914LclRdee8WwWP+xVCsghQTfQLzqv
IXL0ee2esdKgcf2/stBsnrHfFwE+rr+qUffjLTlupGfQOXYjn4l+H6anflREFbPV/bK5Ze9ARkdL
/zoxICIwWG1kptttrhF4G5eXjQFRGQLqM2in7C4RFK+rybNPsM0eReDmaumPJDsHXITRYRWUZLT+
LL2kj3V/8WwfWhm+kpCqK10xze6ohCTR3IGnEwWQVc3tbrHDNvsKcDJ7u4g9TpZGHBJq4wHC6Dfi
F/hb6kMYXh8N3zxJhNbqjzZlN5LLAwBbSltMCM9+cOSNFsga1n3+EgUODcXDSnpkFKUvfUIg5OrN
MzWV9IDAQEa8VRRNVKpn3JfuCNmJpFIfb5YfqcFrxnJg3ABSGbVBHeVY+WX/j3muPQGE8TvKje/J
kOwf8xYk7a3bt2Kw4MynrL2F+9KeEmhVNxl5VyHReokBSQFhhwg29Jp4nhg1p+La6OJrHXFdSgvu
ahKE0GWYV5C+0QdEOMzUdO918ekgp3V3JzeGV11/Kmg+IT/RYbmG4sS3AwpQbtJUKhmVeTF2qr4V
Rn5OIeSfbUPGgsYMvwrXszDPp3oP/4FHXIyvzIs1YaGVUHWgRo+R1UUMrVaFHM+MATF/GkI+xe2a
hIvLQEpMpbyQVIO/exdCrXMn+xAbBbSXZ+JrcFGBLPX/Y+wqV+Zzu0mYWalriGm62koSAY/jg45u
bkRcZA+tcAr1nBvWbXaaAPLTvkz9xwgtiO8OuRUV4RF0mheJKStmbxbSrFnQ0ty4q/LxnkFzW7RU
ivAw7MuGtDmOXs+bNucNPP0/Zf0aSHmqd4JHugegiMeimAVxBQ4u2eCXkLs01AwAy5cJj8STVQbO
empj8vwy8bLcvy+2i9J2Iu+JlkbW1v1yvGSPFPmN8/9KFDXyOO0h6kAJiPQcO6xQgIhHXRWeuoYz
KeuIy75LRnMA9W1q/ECAQoLMPdFF2O+woASGfvDifAe1Wlrnt2ck3PgnM5lBWfuUMpNSoW87td95
87mIMpgGptve0U9Hac9FtQdZD4FIJwo6rn/rasP75/WVRZ/6o9IYMQ7FpeYI6EHo0MLKupa2NPZb
iY3CTLlbgzosVCZ06frNNuYiGNM7c92W8wPSpiSXVuTX0ixMAz3qaI/7HUtLpJyfk6MXWytehplT
JEgx/fqzyRYdleEF2hOQoPo81R+V7sTMxI+CykOKH4l2pGasTIhnP5imDBODO3h2Enu+6w7ZoHa1
LMpqUULJuoU84MBtUvkif+C/AB7lAaG231T7s6QDrLRz/853HULgu/foC/Hy2X7EF0WKqyxHN2tA
yfjwjcGT22dBbcEyyA6Dz6k8T4PqEPcdcYmbUprwn5eyvPCq/CZRIgOIKyw3+yn//IMkuKvuyqhz
dy1xNtTTL0k38c1lDKdr6mK9K3oZIQQsDexN4BZ+HikpzYSfOsihVRpnfqxk4YeB1uE3lMJaBmP/
FwQtWtAhwg+i/X0GxqrsBhsNWU7K/Eq10vZTd9PQ5oAUjbc6f0tUtcSQ56Z2tRKpw1+8OQmd6n4O
7UQgfxB5HgO7DbyK5g3d7RPqI8kEyjbD+itvZEdf/v57FqaaLnGBf5QlN06L0ScMSPZBWp4l9Itj
P59NLKhZYfVQoTdYQOcgu0uavnsuPyuhawDYo1vGJUciDzCSzuV7yQKKR0/2xgR04hgBLMICoIpD
nY+opx4Z/nxF8XbvNvBZXVTXX0Ob2RbYRK5AjHtjYCr7ziulBLAFGlNziF5OoapEH8kPLRUYbY5Y
QlQqNisH5mdG185FFDnTv4b27n49VcRaRT650aAmihoMTIz2EVUNUuSlOVZMILqWOCKx+fjlB93Z
QBHGB0vu35A1I3mXMh2sM0tUbbK5BYjSYA5KTEOEVtSQzva+kz3GeciIkGQgSR8MILfDN0tFQCYY
sNuIlpzcamBueQ27p8lvAuVWfxNqWQVZjCxey+Rk19lor7Siltfg089gBUzQtd0nKCV+spJXbJr8
xC5BsfjFbq1Z9lLNfR4NKQkbvnW7yrd+3zoEdt7bBS2vjCodZgGeaXTWkWoE8buZmo3TI/d//2qW
VV34xJ06iBQEyy6EBWg0or+/YtmCNwY8xfO3egOmbmgkKH/+sGOidibdOkXnKdi73kvDRxpkePmt
0ATvL/Yz4Hw58KIurv6Tfq6u7QoEu1hMnB0U0z0TLgcDPyjLZkF6G349ku9Jg8IXg6QNnte9JPNo
/52QiQMttRxpJXJ5lRGGLSO0XJMZL3yPQAhGoHnYLnwZdsN7iYi9UvKYCazZ4QmBpyDuZ6s6f1+h
wKhdXLCD8SgkYPjHXcqrIgtNgE4om/+Na0NX3Q7/Fv5loFr16Rw0gEsauPmGgvN+swxHBp22JZ3b
XU9owF46EFn2RuX/G3EcmsOYxkegwkrtlR2r8f6btscelUmqQupProMzEHb/mWCeCs+J6xbAtAaW
IgIOWNHEE5UdHk5Ziaejac32NimZc8UOEhLrNZ15ZfAhz2jjNo4BWaTpGKDwyRr97wAEHwoERcJn
T7geA3Go/22S7nzAHr+C1a4gXA1a6ZxZXRMGlonsM6UJt658StM/TcnJ+3W0Zf45Xxf0YmCVQqvp
6Kr0Ju+jlJEE45Yhl+cM4jinOH+AevRbDbJNMnN838/OmkMyZEfRvYcGNcbkngjDcLgdrjIHYO5V
vYlEjdadVCyAqScnFX9Xby/u6TOaSfG1ALInxMj2e2L+mhkq7mNdWKng7Vsvh/PYA5OyPZAAe4pZ
w3rtc3D32dKJ+Zwck5dsDi3/XOQmlTRZEJd3SONCR3d64aHfiRhVbRJ7I+s20aYkKj3j3hfcX+UR
cNk27EoM+8+X0g7QYwLKw5Ow5d6XKcAreYhcNYzmH5qTSuDObalGeVzbOi6tUQ/K6v7uEVXVkkLD
zlbi67uWEBrp6QHrvIzQl2IRwTfOILIvDR2izPY+NAFyldpToI2QLHnbWTdMF3HNY6Js5Zdbcun6
6cD8qjtZn60C8H4L9OcLU5Iy+6gfCkLkAdrJihjp6uj89rPfV/v57jYti1TpJBM4nrGQ7FE7FWEl
hxdteZchQZjnciySmGB7qwEF+5CIeT5Ln/22rJqgnN5cXNTIqrVzkRTa3ob3pa8GevlMgAo76Lyy
sAKfsQyNOB2ptg/OYwhH+u2FxZGNd2tgeG8OQJGiQW7QUXDvaK5sEmouUxz6wUbldPsR1og4uSRy
+DeXqr7p5V9gpKjrhD9jqzpmZl6QjsPbLLDLMf+oK27kLfh2jLfOqpgf5FR+ElMTfA3X5HmmakVg
uc+6ukWNePk1TL/f1woXU9mKv9KdiSJILSgC0AtC/0F0230lAegfwq2KA6OcMwxRUvrl+g9I8VAx
MWWHmR5tINxVew7PDu3uLXiKADCc33SVyknwn7Xqan8iypfC5HGDW+P6ST/v8XeGdalqX4XqULJ5
a8BsHK1UEvGbvh6BxT9xCtUlZzTXF/ZeVmRzzwHvCWQj1RMcxf+Q8alRjy8y8mix01d7u/753p6c
z4CRgL94OPQhzrSnRefn71dliwRw/tk12U6yKQHo77KaJ4w9rrWTqlQk4dE3ilJiOKDKpjKsNGan
8SW4bVzNyuSNAyDJ/uE10IbQuZB5n0JXg2W+y+4GWS2XHulT5Nwzsk+Aqrvo+sV4u5rTov3wcmqK
JzYALyzgxaVLuedGJRb1F6q4EtixvyOKETSTfzVEglus0ut64RO1OWGzakQVvTZzrNq42/SCuvRj
TaKF7ftWY3Xd2TGPaJHdngBv2d9AaJKw6B4HVW418uvAT47Sv3Ro2aZxt1+w5pY/wdsvTzFLcQo4
yoE9c0Q1uo1kkkvLlEWEgSggD+vcXDA/oPFY2K8f5pZ4cA9s0/Usauqhcqx8ka0LIq7loYNvXuds
SalSRLsqCRhIvwsjgmSo3psdAWD1C7FsQPMg/t0Vad6h1mFebS9wo0ZMnO6E/He9uVaPNazguMVW
KfyfnmaHufvkRhx/pxW1G5RjWg1hDKAtJOu7UrM4oH+csIJnXrQzE1Ra579F0todLfE3INmFzqUJ
9+7tmeJKlxiL5jeuJUdv6Q2YnOBkEcsWxoJUPJsudNVkdvQx2Lbq6c9mHTYz+5asagjYVLikc4CB
lBDvLuJPQa6iYPug9tUtXRgXIq2P6d/7uiMChXUBeA/6S05VGr5gDLD219MzGc0oFT+W6dm+QpxF
XqlWCT044YG2GWJm4jlfYMDb6jRQ9JR8E+PsCeE62KPBy8nM0ts3tBM5kcNvjr5aKtbFKxGiJ1Ol
JTjUflCpaxjfF43H3pmcny6VFoPxrOpCRCQIUpUB4EATFwNsrUmh1MWrCfDo+HRMdv8IlsvRC43x
cbHZTsDvvcvu69iCHzfncoPiGnPVBSmTbu7D/T+ltEHYwlXn8DiilWlgv7Ph0LmXqIPMedpTGMls
NvW3DIDayOP0sW3keJ4xMK4XOQK1rMNaCHIeVM8fGAte75i6hFYMOGN9fJ41Rgp3Y2Jni+bNiDyT
hfg+ZYWXapW/UvnG3Rid/zGWuio1sgiK4po2GuD4vMs/XVVmHGCjHYsWV7EpoN4rtfFctZOq0cLH
u2oLv9Cdz1uYMX9IhJ1ekFguq+QdywOpS7iWjTaaQDipI4G8Sa4DQctGUce0mo3eHSixZnMsmjCn
ZqJQcwm8i60r7U2feUJUWqEYerHJrNR2j0UBrW0YM0FZggVGMNsqLEqgfhUtwRHuOqwvzC4XyqKP
nKHWA00vC7iGpLU/ALPghBEiReFZL3FOhBscuaGtHqgK12+Aeeu9LtiP3F7msiHzcLAZM0/qAky2
hZ5XGzBmPaQoz9hgv/QQbsS0cLskQXKyBXK5egULrXWxOa6Au5TJcqkKQY8wrLIn7WIXA7PPf8Im
L86SGeqRE6lRslrpJ2CViAdD8N4knpEoEYcDk0URZlkj7tz2pAw8ZvGXGRhpdK/BW/Nn2NFpQzRE
5JLtgTaqJmYTx3T7SjWstajB+FX367Ema/Ktm3UwvBXpxADAD9YBa4tpi7K4ahD3cgldMbrWForI
Er5ovuAC1JzyTzghu1nJWq8aO7mEP/HznPRyKb4u3UvwyigG6uPUQZcevLYu76yinuVrBJjQQi60
fN3R6Xvzrg7mnYrYa65guqqsTvkkZMldvaZqOPMqtWHCIjrwd/T6maw5Un9Ano5hs06zhtzxaQJU
cXRZhJhl/JhwlgP+ECRZG/+OsT/dqc+NHKiMRnpaUUzLWDlraTgppi6k/sTVkCb80eWwCpgYfO//
GzBx8cq8GkAUlK7wGYmj/eOufM6X3W2lqkwGbLx2h29VfKSry+Oqabvef3s9QZuRyGCAHJAZoQCR
FE/e6jEgcKNVMbghGU45mNkqJ4KTUgJb2qmKs0rhN6LX7r86vbD5l2eOvM1Cgn+4K1P00tctGR3O
F/pyc8m9qm7KpikMO1xyiTP1daWrBe+KoGFVUnc9/+9D8mYMRav24n3wf9y8Pz6cYuxi8eZB1iom
ISU9InUjGXYzv0L9fFyDLM4AWRTDBoKPinXCaYZZKTtO4pfVR36d9nuTpUEfKBpAvc9Tbu99srQf
b8Qui4Pl3ABZ2wKjsWgQRVbJtlz7G416oKZ0hczHsp4CzQdZFrmcTrAKGihWXtdSw+UJS70w/b9Z
yk7gGqrizkHGUxn4eW63ZqBVwXAfFZ/JG/SQUVSI5FVjfQxvLnvGogQfYA9/Xf/A7MfmzZavVfjm
P+wP3qz6DRiSccqOVRvBw4ThNQRAZrHHCp0np1JelHc54IPmLQN7ybJqxOmRtpqoT68CG4fSpsC6
ZFjFE7uqZt0zVwr56hYyJ2mESq841quUhqbL2CUpyCBBe8Ace2K6KbKbJM+vlX0lDqpQNR+11BTQ
4Sx4RSDaAmp6ZU4SfL1Et8wlqFwNdrSzI5ZSAP4LCz1iUuIHvwJfNzZxuWh7BlnOUQRrsSQdPK7M
ADyvGN6Eu2YqnmjTQTeSW+vi2D3CkI790jC+0d3Dk7jf/Q1QLGMMGo96NTnclDMZWVAs8j0R6I0s
4EPnfujDvSxVXRD9/zEgGt/j4/SogltGUQWd7+BKRgctCW6qPM0tfttTqjW8x9QQOMpKH3C2vuG9
GWux0rggnWrdGDHDZL9gHAyC74DyUPvSfuewT5mLSN7KjeNScyyJc/iGqyl+jy5Dn8zqXGvtcu8q
QTPSIYk5q7I4iWrNlOUTEk7xPVgBApllG/YJdGiDesZGyI+C8gNpHabcimoRpRlQuBavAcW/iIt+
D9TPoPQi23SidY9pnoeo0IkQbsZyLkPxa4ehGDv+jI+iJliF6GtvW9XPoIiyMLepTTB9WBpjwM0L
bR5/a/z/YhoT9suQ7vGlaNOKMws1xoQdbz4uW96p3KQbkqlBLWC7yWjnBSLQf7zc6QSFP0iZs02M
haejpB6NE37pcqOpPFU+iW3fC8E8LJBolthSHm2va2bBRtw3oq7H0hVG/nINKxGeSp3NJkLFzh5x
Pl6rWqdnbqltZHJAvgjqqhQRXHU7NihmOS3s8PvIeF3V3c1G/f/IEYz5LY+ONKQt1biB1vvoi6vP
c8DTpmBxrWpZAMql/owc/DoNvZSyg3IeEsBN3ufMIibMvxqaa99CeqQJQZLKGogeRLJffC0eHYt+
KVHICvid6WhsqJpdnetGsFGQ7AUC6duG40wnAPdmTcBZuEG1Ap0AxV3nVEYQP2ms0awzNXxHIFqj
OoOdLg2Q6WmsMyOZAFm+5uLMteZEtFg1Mub3IE/5WgLgIZe3RBKKrxD8nRTMA8UgvYNbO/32f6FJ
nUFKcqrGKn9eI+NNcjL5mmm0McAGMmxBDv4wIPB2fQL/Cv9VooD5vexR9WlAD6npD2xxY0BWxQJ+
5aZ2W1KJWXSdRjjHiU/qXfTqDdyM8oYSmbfzn88haHpuYkWX8GXgy6RHqy5JpAkYkjO5bYHduMLF
uBtzSsXQLZ4Uo8au/ELPp9Gai/cH8LHcdBIcuxmD3ckQaWE2jDAFzkd+pPBOKbkfyp3Ea3qCGJum
vr4134MhgMc4LZbqG2eEc/VqG0vE8S13b8/izAmShjwTyERnHFCNM53YYmlhthd0UKieSHv0Th1I
EnSMHgrcjjEjPOLOg/vePQfy5KGtfATks2tW5fEM5y7miLPIiOolybOBl5Ve5vdyrZXpOHKsS819
GcOSgfwvefvANtBLzNYI9hrk7iMGirHLVuSw4kTW03Y8XbWECLaNagM88ZQFiwOzDYRh51AyGQ4O
oGKNmCKUDwBbmAxybXcyaTTFEAr6e2ABnn4GmAyZtahJm6MhmvJu2tCUm6MuAo4kp1K0n2xCiuNS
kg1FrPpUM7dSk1Y4GEW0OpKAeen39d9UKNW6HMC5d0AbXMtncopV6DJqx/gKcj2bwA1O39CUH3wq
Vo1P5LsM61+FZj/7hCbp7drENQq8MBUHJZtp/Y/2lFcf2c9gwgVamD/PGJdONnqafUFRDvn8hBY7
7PLggsNgpR1Ybw3xn9SRzZS/eVpDo/F37VpeTELvEwVTV2x4vtWAEcJz4PABYQ8TjpeL/C99G4d4
7lDu2Ge3sEurWYcxJEOErjMiar9w6TRwuqWEj27Y88MiW7/X7AZDkH098zqCghMVG1dm9kBW3ITZ
YhYtQhl7UrwNhUkJuhR40h9js3LFf/8xkM88kV9AGbuhBtLw/2V3WcBs5bWkaacx7GRLLQD/van3
LmAd8qCDHmoI7EotgejizsENnA4jRiB8e5Fss+FDnAm0TFl0FFj4IMm1WtBpnK9jYWJFn+C5q1+L
Pkzb2aO6EYCzHCJLmbgQatHEBNxCzFQcQKIhJSCgyP4zlFLjTLh+p4ZHNtZdU4yEh99hYek++aF3
8AMyj9JOz3YRA6DxPaCMJudBZFFFQKqwhk/GYV+UFDaxRyIxHoErMA//mx9E2g0gbE1O9Z4ZPpEa
F0qSWjhVoFAJpYHNhAGFrmS1WZM2k1MEmhfJxGckVwxE6UwUQRCWMKBogyNbzqJKXHMQJatj3du2
8XbXXENQoHj386YqUhLcyB/a4Zk0ta/LUBd+8ehalxOemmRSpXGdU6E4G/t+IKN9ZEsUL2uz8pye
NqGBmIfwWNWwrg155jqWudDuulF/fAC3vjiY2faCvDOF87N2abapHs5ieYacfxFr0xU14qz6PHxJ
NAsHYDODB9I0PKbOktiVcJuIRX7wORKQZoDvEkt3dXTZIymgx4/vJnhRSawS2KHk4AsFI4mVYqW5
8CuW8YoonOzhvi+Qi1GFVA+KFwvXHqdAi39qYI6XF02yM0roysflFd6QhimWxGOMKCYnVoLzuGJq
jK30yT69VbUUoqNtkWvMC4BeEQPSGfI4HbePFfL/9V4cLtZOjmF/y4fXIyUbpehe7HvfLhy93fyv
Ew/6uAKQZD0QGiMvNtxJQSVT1fJN4ihLIOuYjMjfRH2rc9a6tW1Gbs5P/jA5VMN5ZzI8UM1BWFId
KsEBT/s0jMJAVrwlURUzIgWjCtGsKR5SgSeM5rP4q0dgaRF4LcBPr2+cFZewNvVLRDIf2HvzJUKS
mBaLT3ieIhJN0bhMJkiOTSabQH9GVza5oOf6V9/sRdsMvA0n5iSaL/q34H+ggsx/MLsRUfKGM0Sk
MjbnF1y9ZxUQ/wyZ16+9i/MK1nzk0udizOQ9J9CaW9pGr0NMeuh4Tp3ijtHsYB/MAGxWVIl9HlsP
03FDR1hUL0i5J4KkkfP6FQCHuTSHVGRzXxt0o01hSaESZgMss7dR95A4s7jgK4oiRA6xiAk2id/Z
DFZChKmai6VcYL4+avE31i1n5flc8Iau2O9UrxT6gTfOCv/x/+tnEs9cHjWcsQmVUnpqvSJs/7d0
6SoIjo+BbR41dGDMUOdl1NHM9WU/yLc10rCaUWzubESpfzuDpK6hICc89ImNozV1LfdWvf1xhcX8
NjRvh89fozBI1eVhu6KQIJevNLVDqnT9aHWXo6VdgxytKKRiUNce5T0ucYKQQq5VS8FXLSrpeS2F
apCe2BNHyawgE20UkTQleQ46yFj7n4rWtiev7oBKeD7uUa2JiI3lTQ6Ek80DVU6DMMqKXnjUZvuV
HFYNpvphGBkjz+RUElwcP/03jValGn2VUQDjaiYOxfZUZw0srvraNjpriDGH9Moo/jR27pWfgRKf
U1g3M0RrVVPgmslEv2fNuRG3cSyZD7qx44A7TV1RzrROe/EqdjUbmkb1uBuDO9zsgQgrfjXDjwjG
SgH3GRzEVsS8NTodRnB0DlFLu7pHg48eQPUYCfDeWW3MQ/SfHen62IhENlv/iHuQTI8wZOBmRDW4
8unx57r2G8QTQtSzKTgbHhld1Nvp9WnCRDc8RnJPZeEFrFDmsmbTcie8Bjsd2GPLMMYmm0VEX3XI
Lkzvwyn+jg4ICVrWHxP6RPh5nCl6SbLvs98vtoEqVRKrVJVjVH8pDK3MhYWCBxUpBAZHN2U2fN77
yjQA87zP4Ycv1A33BIpyGPrV6hkXcQJf6snfJcExGT+Xv1H4X4BqzsO5e/izOtowHiiHPDRQoMae
gzdqY23TcRsngQtrqi+PqL8Tp5HpgHi4sTQTQ5dRgNjqmynuXONIWtJxPX5Mc/1utLMrtBjN0W7g
d9HyFAq/i62HWR2M3kAdL8ZgMW1NP3Dn3+z0Pf2ArGCB0xxr82hN0LMybk1uKuJgUS4546gCWdRs
5pIbPVjE1W1f3TcsYJrwx60mdGfCCQJrHIDfqLbfktAgR0lA+LAGRYhmUuu9/o58HOVsnwItyZ+Y
umYOdS/dTgkbT1IShEG4pEkDLpX96F45VoRWbaJtmA2xCQcRYyvz0F7EuTNLQTYkPSI8FdYJUqCB
PrK2+tuTvFTA8g6DojDPYFeafX3DEHebVM+EJ15cF+I58Dvb1/mMgJUNDkcQ/TvTF5YHrWHh+DpT
6PSiL5DQ5ye1+cRF8lzWRn6bWnQKeWpeprzqH7/hgNmvq8d80UZ8XGPSMaKwk0mTdEO6W2Fy+xO8
4B7Ezg8pmDO4jgtnO5KNKOwW1qa26uRtSLHWYiwSMCJEXG9qhs+jvVUFWKayXiLKPGlMX/Or0/Kn
578XrwgDSda81CwAXxI5EjdGFjdbuL+CulQd2Va6Zc+3qcHyASmNb04k1WEahgxpuwsB8HRnIJfr
ZC7sFzaoK70o+yF/iG24j7ss9fBJ2tZuiyInkzjsHtXwHlsXv9NSkBfQvP//kRHoGP52XA6j7Dyq
Ds6Wszk4AWeXG2l/Y6TraK7Z5QnKIFasAYk3CJckgYH0SF2VKXQESv6BAUvhUGOhRQx2Pq9hk5kg
AGHsuYR2DAq5QrIJXP7x8NySRdeROGVe/DdFvBC57n5MZTZSX5K9LmcQprKFm9MR1xUbdfsJxCaL
13nod9rousz2NQ76dCG/TS6PyNu1BMQdlR6ZKeUa+B3g6PNlXmInr7EjIDU78/s1WH8bgA28zHJD
Z2pcFrHiygJLYJsrh7NUV9RPlPqpDRlj1uORszz6wJH5AyW/zDQGTFfoLcP1vrW/Ay9HHyZIO26w
VB2VRbyp1GIhY88jt9yjl+fFrWHoXv1GUg3uNYRSD3RgpuoIV1lUNskQIzuCgjbpL4qLX8cllBm3
H685cVMGQpCcrzEcVNOfmvqD7zXI8sHUoUsO7auZ/L8guf2qiESWYcPiG52l4/05dAVvm0kFNxoX
51fdiKJiY0KBcH/PsxBz+WVEvyo/DgZmm/9bR/6hqFLXd3H1F1xMe1BVSbz0ywDrZw9tJt5lhV4O
aXkakiBy4+a/r0SWnj5s9X44Q47+3eP/HAURDQWfXeEBFl+VoaD/XmZRph+nPyIcNXWtJRvYAoPh
lSNLvRzi+Pqef4kECFLKPmlJlVoNUBAzyYsY6nLSm912EeAAfq2WuI117nbbTMnDZ2qSTF4ChHV5
zfcNPbqL40+KH45hxQjKWQAJTkBJdmU0ZHh7LHrli82SAaP3RP6BQogtJ4R0A8ok7aYM92ufrlVJ
S6BEgjKxL6OvdBzuHVkmOQ7XjucwbZBdlqkNjpwQnxvoPqvxPht8jNULtP1DhmaGbusqFOLpeSq7
q5BCyz2emHwPrSZkgDihRCIt3lh4D2vXeRkhTfAQUdxF5xSIjmgTW8t9ZVLnzjZHgFFJNMSbundY
K5j9QMYg6eUBDm5Ql7ms2YcIkw8UccYJRW7uPEOmdukUUuw5AUmBk7gZ5TjL+M6kiZ9xTNAQzjXT
DqSp5ifpgCoWpqo2EOfBcaENwXkzt4qSTG2eZKQx+TylvCnO6seT6BQD8TDjYll3NbW1j31HtNf+
KVfOSOz5BQ0UrD+SXAlwtI3QwWkqAkhZTfTlcxaq3KgiOnJGtWc4gmsVTfSjFj9YqakRiZGt0/tx
rWDfRiud93u0lFYBJsqf0k/uO0fxY7FGywtWV/KpnUUz06yT3lgj+CeqLl1ceT1EQMtR8i8t6hhX
vLv0csiQZSHI+4Av130aW5CfiQ8H79Uy+ZDcv4uT+e0/dcg01I0XpsOmPXElV7Ou/ntNcXg1hJ+w
ok11BhehDvgv3ytRtd7/7xUNhZ6AVQ45tofJlWMyK02sXv/k1hwkXuV6vaooIvN9q08EmsH5uyK5
PF4ENX8xEuAOv94RH3HdUZsBVn55hCM+TXWeeh6sN300+ezregT8hj4x3rQj8u/NsZV3CPAneoOG
K/AP5C/ZoioG5kaYoIrdtm32278wTE6S+zLUwTN7/GwYy+pcl9aqCvsLKaKbJBsLXcvHDM13OCfv
M/TcFc0Lj28EaN2uPw0wfdPf8vZnzvPR64ZT3PQbtJVNvB4D2mu04mkmjr3w/9nh5rSFeK9DSooq
9tvJJgUoXZrz8yObeiA8s/IOFQKxdxf2oQMS82D4nC2fNA2dPBPGFAOAKOcVyHTy0yinECJsQX6R
m73GD8eDRfSZQs3q6fZf/xnrlLCJaB5bX/E9/hrw4vArjJl1vsLjueWK8Bl30FAxZoDCtdA3Ju9u
eadxNuSDTUU+iniI9gSr4PBFBWAZ86esDadvVl7vpz6O31UFSca14gTVxojqar0Tvlu357k0V2Jv
FREsYRXSkPx1gTKwEeN1jR/3wQcrHTjUChaS2jKB4sRecslGVH5y71/toD4+P78YDU+vtOXKuf/J
4NiyqJVzOz+klhMuKjlwnSIFkn0DoRVImOnokssDfcqdfUzQ6bflm7H0FO2lnHC7QswEvDLAbsk1
mlGhbxOjUWVvzeOY7IZ9F8LbnNiNis4W5b1EMaM1oVSp7LNqTU2ah0zJ3XAnk5icR5mrrqIGCL/M
3nlPcBRHRrqjZJsL/2vWg3Tj9PuIW5aTdogsiuTAX9gtV1XGgVlFkQdhDiD7tz/Y0jnwVxMp6nhu
veQlsdPlLWtDk5v/xfVyvUIn2TfIGamz/MySRAGhW9VVppOJb6bMZzXKfpURXi4ZkNkPEZjaNtcs
S31s6lQvZSA7qnbrJ/uUjasJiu36nOPikD4T54EjSVmbaXcFnek5TWXq6AUEYPgruh+O4oTM6L2z
9JA8/zVvdBfteWbsolj9g+W6+eJx5JkbrU/wy+O5M13sd69uiRrK5IaQ2NR8K2YCQvW0NlnEBvli
W3b/HLbRPzHmmibO+ygi3IRmbuS1ZrwsGwZkJnBlI3i1zwz3knvQHTOq9tyzNl3Dc7EGEcMmO9Sd
wXBPI89QeTHPyCqlLBq9wrJp0UsBdk4z7GFzwx0F7LtbI6sBqv37Ba+C79bafFyzgfBiaRrW4KaX
OpS1hQ6pHdQJ3CuUZtyRx4EnI/PbahdnPsE2cvBBe5t+6sFUaOkBxB5tExkBWbpWiM0KTn0l0Oov
YiHqCbbt5fFe8gOmLFq/qihy517KCsC0nD7hN3pc7khLjeVnnwYP+9SU+4O8Al9a/OpbQm8eYJfO
DQl4TVXAuCrQs1ORdvr1WUYBh9vrtpUz3ZWxkYJe4Bg9S2Wz1Ew4/qwJPB8xiYl9Z6p3HeOKEcDP
1Nyzjf3VODuFHapTPJ1jVhN9rVSVq9AJzr6WVZ2Y0MDwq5VAtvb8+KdCaMQ6rnBIGIueVeFFW3PF
QsMxtndiXKLgjbCclXlICUQqnPN95WYnC9FKlT+G0z2eBLyrRDsz/qRdXsT0p1SPsDkX6HB+CE3i
/1yVS8KrAz9xbZNLiZySVoF3y46Hq/BA3EN15tQmLOM2ZPgyK6fKXr0QDice1Kvg++pLc4LJm/uO
X6s8Q7/TCtMM6hLxouZGG89jW8UE8NLAy0BW10nJHFTn9rwUMqb7EbQgApEbZn2FgtaRoxm2NhKL
eHL0sCA/7/9MUdubD00mntkKOE+DyLGohD97tMl82bWd3ZVutg8xhPmL/H0VaSMFcKBGMQnqyPtl
H5zt4YdT0ifrm00zgqeHhrPW4/dJ4+1l24tNtUi/nJAKToHhbHyupHvn5DWU71MZXGmH8xt+oO+s
Qc51z2LzeHHQ6MFjZLNQOgUKox0e6VrcKpNXGotFgx/XWrqpMhLuFmO+t0Qi9Z0cVjkVCE1dXzlm
e+mCy9dVpNnfH2A6JWDbM2LVTH6ylx3rsFFxpI/LxBl/ZGI1I6bCMnAuvY7jEhjhGgM3Dt8rOiu4
bPJ0QxEGUmoz8pi1dZu3DaCsrpo5sARIqqpY+LT+8rIuT6YwMkZI+35DK4PynxRRkO2K0jG8e0x1
jg5RN+/evy04Ijc2gxL9eQWH9dSkkPs24sKDRlhWbmnfvGX+zOpjNdI4tw8ud8uA8++bUrtuw9u2
7ArMSK5RGBBYPW8QO+sg+5sk8p8gULpkYYVxggTOzNMLYOF7+w6E5GA5OKa5epMvJ0PMzBJnc/ql
MaMb3HBzAHFCPBMgsAs6JuDxb08WdF4mHv9+bgdgkwLNsXMow/N9atPJGCsJeymmhQ2P1I1iynKz
eCvOVRTQWjrAGCm2G7lK0UYBxDR2Bu34MVrC9SCfZK8C2J0OIKfQJbryicuyT1cqYAnMzfPxWpF5
UnwsolvXK1azmKcwgJ7wCUijpHKhem2vHLxZjf0+vj5KF7lj4yQCaO49lyHGDNZ7b49YeIJt3oDS
ZWSnhQhGCiv/uAx5REKQI9wh0jLms4UbXd0RuK1XbUaxxXsqkfNKYHhNY/AY1Z9sHImVcj2GJ0hs
5YbTypCvFRELAzxMi5+EZrupz88NQ4RGed+3tSY5gincphK9PdYY7sfjaM3xY4cAwDNQSNH7f0qw
r1eTEuLgXrk1odmn5xwO34aqflVERY3c0/5jCna+fOf2RveJ4cjYLbTR4EgfthG8PP3j1nfhz4yT
Bt9nacKKjL5CVq78oeN6AHuDuBzM0cGTw4GWpDt+UQ+x7PxACNGXEIRJM0tdr7s0rFk2QaOw7NAk
folhcZ+h2Evpq+n6Vb9NfFfBfIhzEwbDaCxgPT721ttx0/FONt0lA13QBKpEuQtPhoINBVxAIk3X
zVDcKHAilnPC17zwimvCn8ViThRepkd1Z1stlp8vaOG7O5hZ9/EM5GyayvgSjXB+tnaiR+bLnFCw
wy36xpFnWf/kqCg2KFD64EpDN9VEkSAAE/xvkTNbSFGZGoQm8ZbE11xbBY8vs0Lf1rAZU5ZvN8I0
irtNOB1pD1PdfErEltSNyH9Emqv4ne3kfTc1/8AgUPLwKwcZgwgoI5uumFcLsnm0kjhTz3vUZOOa
bxfBazrf7YYPCIk9K5ZMbCvZlNkcxMKJIlcTQPwBdbAf5sdT54qlNY9ztog/fi6UCTnxWzNg0diR
XJdUb/BTmIQDvmEFMilRiU7nDFAVkrcHYnOh6ydkl8Xn49Jzc1pup6Q2SNyNXp/nDhiCi07w8dx6
Vf9UCGWRea3CiGBpmxgXUtRbNmVyLctMoaxYHFzoXEwNt8ZBCn/g0BcJUarWaJPzEuC+558GUBVV
++1+3qBWiA40RrJ98KNpBTW1X3YPOPUULX3zVuhCirQa8OVDsIPhlh3BWfvpKAoAXkFpSCrcSMD1
tNHBpD2/aZeY7WE+BlmqWgrySZxyzlpw5z2vi26/MhrpF4oTc50Q0br2OWgrxomCgib65oeI+Ajm
PLgS91WMkzc+k+2UuiMqENJtx87WAodpTrfeBN5jS3IcYZkOBr+Zi1bI6zznHHhot1eeiNEMX8pA
/N11/Het3TDFyjsOh2PbvAHt3apKujCBS5bcfyw1pZCWJmUafVLKzebWc8SRuIBv7/eFyTAPo0k+
HUZtLyBFdgh7tUdYkb4iq4NCQ81PzhJ73OZfdX3fD+6lXYTOXD+NVLBbfViAOYJTIKYNgG2o1Qs8
v+LVMM+cEphLKJjJoEnEsrB/1axmRIAaWfTeE6EMy5be32vPnIC09S12gdFT1lOOVXo6OEdSLFU0
Af6va96LqaqNE92ek2dgqXxVNlr5h6rHsH15LWbl36X6EbUW5aLAW9dVgftmOh9Py3v1cygJk8F4
9Y/sPrLzUsJ5ztrlNWhJaGXSTfuoxxt6f5zD3wLzHMtgqPiv64xffTmLbXP/bz5WlR0r2qUexrwE
5Q+kXz1KC56eQbgcoKhBSJQFDcrbQajyLiHkZBBPL5UcWwv5nmfrjgq+DWSVCSlATZNIiDJeTBaP
t65zQeD/XlUOtxyJdiy9XCRVY2ivcBw5BWXZMRLixVjgOsjsKKzGH+aUfwc2ZQfQeu9t76fAc+Bh
RXkzabTM/lmLkgLIOXN1i2J77WEebROL9sDHZ2h5O0aJlbJkpS3MNnldgnPvJU2tUSyqZvuXM9Am
TIgWBhXYLi11KcS7xSDVgTVO5ca+HqDF3j6tcAz24QWZ2CzFw3SsXCTbp5yMnduJ0tbi8UwD7ErK
d0TRrWmvgoFO9gAOAy/b76BCAQs5yqsqc1mAjEunOZDYWGGhduYxIp059SrIcXzNvwirjARPmDrD
WlKI+XsYhhNdakM+5ra+JavYh2Op/Up5Dow1/ZM2iaLNT+QZ0QVYJH5PwBJwCFLMZSxjoBCQsv6u
5VNWerDfLD6YgdFOCmF1qbn0fe1Zo3O6GDp01IxAHA9gY26a6VLWG5iBpNCqhEOh4j3Hfn/R0EBJ
kbAbiHeYgwKuKqGV6e3pceLH1w3dH576dvW6qzpC1kUm+3NM9n9k+ZDynVhsY1xprSFyRyRDmjO7
HWjIT0IyxPhTqQe0phBr5v/Q2qG4TNd1EW8sPbuuIAc1EITsdKCkWmBa/55GfItCpSzEYyYcrrHo
Z9bhvWtAp/hyUJgTMYcm04VQlG9qeGjWViLKxkYXAY4ZBh/EKy6zdH9kzVkTtUXR7Lx+FGoE7t3o
qrxH9g8SSmU4EoNJksinPihrl79GB+EQspJzOjv2NRLk0dJEfR7AE6fcOBRk+upCbxW1Ynq68Lxk
RmhmuzB0zNAMazyGqH+t7cugYA7jXx/zPPx6CB27KNU7Phm5yuth7HT2BdcSHysL4QjRJkB3M/Ob
xecGTfzDxYrXSC2YAQzZAvK/8qiMp8G591X+ShpqFXagjVzt7oR3RGvJ3kYekOLycRzatLEf39Uu
pJQJPr5bn94hvJlonKdNylhRxYOYDX2Xq78DvdnNwR3LOE+g1flQ7+86gYMq4JBteF2PTp1A0Fgu
O/XJegYwB+0yxiao3W1CVOV79fHWQP3+mEAOJy4fxXI8Oee+uIXwclCXLG7Pmq+ZNGEgbT4inDZ4
lpr4rmVMmalgJdJQ6gALKIFvPisrmQiw7clevoCygxZmnDcsiOhIZAJhogwpi6A1wdJC7fUwmYZZ
4dyGJQ3MUepc3NvvnrpMhR7oWlWE3YjOeBUfdkD3Eiz9mecjBjeEWw/G2nTN7+z322dk9j4MTz0V
9jsMLX6ZqUhP7LjMRb6z3Fjv18XAMsMkLIUQXz9FjUJg53RGjRWvnBsT7hq3BpJF4KOYRW4oayLK
VVXkrSnd8R4QNeQCzya7gmFtyreQlDQYCDfj7cRTTRBGL7pDGaKW3P9kVg8t/tsFyeXZNHKTAj+b
gdD6ivtulSymdg/tApwDG3v9sOeqNf8dMUj4ny0F1WLEvkfpBx9Y83gGRRS94pjkAO3camZXXouA
H2tO+h1+iE0Tge1thn1W1xQxjqQWgEL8EMyRRHiFUdU8rO9/LTAY/haQBDy14Ps4/4IQlkkKYrQe
nJ81nCmx/tg6697D5cHFYVV9eXmbs8LZnHVIRMY0QU/eUoxUvpGLmEXrkcmj9bKZrnBoNmE1vzdN
g51O8HM2Nb8k411VQI+QMwze7FBkodXiAKXk9pBvyt1WSgh3beDCOIVcp5Fpo+feg/qDuWZMy4cy
D0swe96LseG8mZIW3jL/7gppSfZqUcnejPtl8AxzOCSt8Zm1hcUbXxASMUVn3k04whBkwfRzfUnN
RuselDNOwRVYPQS5zf1CHHtsfvRJwTvPZi+et57Im7HyIckosgcNGp+kDe6IyOlDm4yIDj2vCalP
zEhfFZEtx3EVG3+9Gu0VniozramkRDfP1oEphTeb7pYEdzUgcyu3snTXwAs5nchEO/vZen4nipqG
nDtBfrM0ujvc+Yv1JwyfyHsbqsshYJwTZcCgWU8wPOt9for6y/tqMqELcqzqEfD0ch1BnIbSjLWr
+8Dn1Hm38huhRWuX+G8heDZSDkUWVXS8OaYqQJyZUB/+2YSF/Nd7/WW7CFhCTaUcCpWKGz6kUeDO
arrLirQTfdmpls1YdcGQhb477AefHBIGgcYU+yKi8okB9cV3kUYRzuX7YcaXnMYmCeAuNoxLokVo
IUEbbLCuX5HkbsFF4PxzkqYSGbYLP7nWryHBsgLTri84OQS8F4egmGEy968wdlUAOx3hRH2DR3qe
c19xBxjTKzbDttz047TcyFgQ99Ojt8Z4nDe28pKbJImxgdI4DRMbtrJsDvIIJmZg1XKKTHrFYACl
e7k8B8Yn2eP2Y7mwffLZ5xHR2splKZf3EgMwLHWL6+a+DDZxBsa3HaDJEDhZ6P68xM5xcGbDgURh
f0HMFDbfYocLpynhXRYMnJI5zOfe4dZWxVCswJJngBB0hTbYzbrmGVd7ie9sogeRMJ1I45fruzAw
D2/P/fQXWG2TDq7xEJ02Fu2y07wMub2YYtRD3znpF+MQr0KtpnQ6loAT+5J2VqxRA3tMTa/jFXR9
GZcWBBc18XErYdU7qnzUNDqwqbWkilnoS5xeRc0H0kAVE/Gu+X0OWEuTWv0x8c5rK+dyh2BdVwYK
OITp6dzbN8A3WN/AAO/SKytKoKfBFrpyoEugvKUc4fkfX8Kuz5x3zJ60Usmo0dRvq5NgrVX1Y1Bz
u7I6oX7l1CD3af8qyKhs9RDoF6TYukP2LG1O+OiJE3iybrRGqL+uQQhD+rbvjpF/T45nGUDzZNXw
gOAislGJ58odQWE0JLNdOgY4w66qbz7AuqNDk5/JUJu9INJposUmiGB/ixWNfpaozyK0MG8dDTsS
B463lPDVRvpUUW+nyqV33t9udOEgg6sdJHUuf9gN9mpB31YWK6CRRhMpz/xSFyeyuw6wK449HaC2
B38FV1mHABleyCFMWDSmYIhwmKtfR7ZTtsa6QC9WjG0mc35vIAOqbY/Ekezfals2T+c0Cd/Y/1Z+
YbA1DqOGz1zCkByf4muR4lj5r5GHTbhcGvVeKSbYNMoxoy5KciTRW5tx9Fo+26kzV6V0iC3s4Y0v
yqKpy6d+XE2/m0SxaCWcNrc1qTxWLlBLqT5yK18yIOHFuh2ma9s1sb9BuOBzdQOGcBe+hQc1PddM
MdbKht6VSPKs0Z4KpC1fjEsAXkS5434JqgfqoUxN1uPaRaYf+orOF45HhFBYV3z04rG+QkWOXHdH
BtKJM/rAn7hkC9kzwi13dem6wGHwGSXBXeJRaqU5MATDYlXTnZa08iZVsT9Mnt4vubtHzvPrOU6b
NuURFOcLNnEvx9DAzhvCx3q8oyGR/HtdGLv7WAQlio4Gmnh1bvyJnu3/4D+yPlyl8klBNd+lgKds
f3APddnSrFBUqFcvslyM2yEM9TVUJUl+ExD+AoZJPYluVm1vjBeMmWDbDu0+8ioLYp1BY38tXjTB
0pDGrukB0vpkHspQ0UY02asfCXuIeRhXnksauQLjArR8GknHg22pn7/NqGnTHzqhjTs5gNLzct2c
uW0H20tHpmXHTL0ibMImRGF1k37Xlh81taODTkqERrIv29Q/VwKn84EyUV5eC5OPT921dI2Rds3e
RevQ0QvNLlSSiTTlDpCxNi3hbWmU+IWwRD8bo8zc4S2yS2niobCF3BLsJDlTvAEWk8RNpgu3dj8A
vIjupQMeak2rNJrxXFJ9mFg+P1e5KK2pIEBDTWNeZe96yIqCDIqGKQIKwdoRTloJeJUcRo65paI6
OgFhtkSAy5caTFVhp8/rEE1z1KBJqSF1HAbOq08ObkgTPGe2VbS4qSgkgl4mKEZN60RUjn1WaD57
leJt0Xf8/muP4nsg7U2MYVgSFm+oJlro+ICqpauXjqcMJv14fpPPwzaeKBErdmuTGcrtKoFBSyo2
ij6oC/iZvqzOpHxkMlWjVDFtaFP5kdhzdiNRIl+v8pHkFzknri6fYMaBsDhyKd9hTy9etAdNdsd6
DVaE/GmHmTnxz+ghrALwEmqEBG/tN/IVoqzCsEIZfEO3nUREq6aY0V/4xveMRHgyJTHTiXmQ5NIT
xe2fUgA5ZLsimRelmgfi0PpKDpuOPpnhfeLmfYc3jcCCznPSp+JA2DNZCs5IUkpmQdqXsh0SFYT5
7vB8N1lZ+jYFg9Tq55u4rNCFAl+3Z2qT412ufq7Sh1AuCYhiG7aZP2JNX/oBKNmV+00HDY7bpB6C
fovNlm4mgN2GXFhDEowlSioiQ2DIeRIh9lYC7azmyrMKgZRGzxwIXT72aH1XYM1Zxkm2wXbwSMsc
itSwXq6/C0ZetcTR5vVqajSpvONOJZEp88JfPy4KJbtuCII/L1JEk53ThGdrT1o9aMM4fJ4OB6As
R8s3e2iFz/kjdkzo0XEV1p029X515ayfMHbkw++lmUxz3dOO7oOipSiwqcOpZ1tNUcimao+SBQpD
UgiXZ3BJ6XTXdfFstifIaG09mNVF4jIEPQnmWsuAa1UEv8NewhlaPc+7Fdfk4heppw0ukrGYolf8
dpfR1yF5Q0TnSXSk9otXZ6fxBuOKbZNt4775GJ8F9Paf+hcYXsmpYR4+/qxD6RJPZPsIW8jGXhge
7HOwJ6qEJEf5Uw+HLdAkCHx0zMSSD0KkOcZwQbHgzei4Nu5yoiFOz9+fRucosapmT5ssBM9+VgMb
SIX42FIlB6ghGnF56iVC+v07hD8aijTyKN0Dt5QKJk0Mcto40Gv0HEicjhSwq4c6jx5t3VSXUCxM
zTvFCxXyXZz4rxWb1IBGqkLb2ECkKhhZ0AZk1MowbSEHa7tRAlT7e+R1AP6MGoSsGxd0DxUn2d4s
aBUbRvW2CtiwlFrnnjOvcNrd9zFBl2DwOVF9s1+gIMhRhuc6+dw0bHUcTixggQzPNe0FwigDMhAv
MZ20B4k9UL3UGCQmEplsOruHO2tWCghMckXmcNj4uyoWg60eVUXlXJSbTop9Ta2RI0a8X/wKHkB6
EaowBIqglUly/I/6PRMMBN2Ko0b6ZOpojPrpoRyLBUwOzRo2kVuGpnj6ItlC78ATC7gUTDnlF7OY
lKHrcwbCUrmEXe8STDu4eER61L7/Ixhr3T+AwC9Edvmu+lrr/iHBNez1JOYRQiE5uqh02LkiAq0n
JztsANSixQNBS9yRv3finuNQszKJnWzJNfY/8SRnq7wQMFmO4fNzVm98si8rF5q56b4QT+RN/XTk
+d2AZ0EGqSSUWJKaU/5fZZnyknOJMOO7ycy8FaGt2jRrSA+SkFoCA5ipLYtPSMMf5EorAnj5hHfH
s9TnU2lQwz18I9EVHqL8OKivxq/mnSsqMk/65T9PAW/nHuxAPKNLMjEAmDnbROBCiDWaU2CuA7dE
cD5lns11Cj4hiic3mIm3Iu+5O2NJNuq1ltinIi1+j3PfQCgGEpAkTMIabx/WkNrQCONSdxAZvgUU
DLcs13oSgQDJGe1qxGyn+26aYNvL9tcMpOHzVO5qhsS6ADzYlH+/bUfT3fOBRvYP/xJjTNkIGOyd
JyqRsgibb/OMzzeepFFXf6XVBKP6c8gXxyxhNagVGpJzkhY1oTCaNFh9bJjzUj02fGcTONUDr9K3
Sku6+VV/zZ4kXdMStCQkUW6xrpBvvKdvURMy73e4QHAGVBL2bb+QutPfj/doaq/AsRstPlgVye3m
g1tUi1nYab9R5c73nsLBx5MXXMNwh/HlB7guoINx5Yiys8cc63OQGumlK6u6c9cHYNTVysS7GGq6
xl6ItGI0FqdWds1qa5TREFG+JUUQSSUMx1gTPzPz4NlmGJ64S7o3ipbvMCU9dda9GU+OPbSCUpWx
43/ZtLEgedy4/WTpsp6zMtcor+2MWTtV9YQN7i0J3FvgpMvNy8eR1VIJwGcx2fG+/hBrgM1T3aVM
bqUaTGUIv+e5dSkFLVEX+QKzCbbzyUJQ5Ys+XBwMMAB+DNlM081YuoTQl9Ju/9lB69eOlrSPYd5g
eI1KuDaVeUOHNJtmNhLh1BeYMqNpJ6Lff3YM0XoJAhP6eAqn2MBsgMAMjoh24TQSeAvZXaKCIcX3
BHN5seF6F1melNlkHA78IG+IFu4Bp3D5MvtZO3Zv8BSxbojqX8uK7gukN8JoQANEzQThwM0hS16u
1m/vMfAHmLRjvwunaWSp0ldbXUqEQj4BSEdfT24VNEdOXtMnGUFP4lUrQ1oyVLummVgr4RIzYhfN
hiUjgXYKUzbeQlJv7uczutrzdDBIW324tJ/6Fhf+XPXU9U2f6s4k744uEhr7nGIXK/5HdRb1OT1g
+u0zkQ5ZO4w1JTB4ThHdW1w3tKvPQmh+kHWSNxPOEeRlqcKJ2U00UWHB7CMd+7X/myvtQhER7ZAG
WBu+wbM2a6ux5ifPF73jKSxVeaOMtOVLpyFXLNxJagYuhU4ohNn5eK4KjafFp3Nn1/KMrPU0cDo0
0jXx8dwC+4JZKNN3+0QeO37cQnBQDx+fBF/td2/wyb/CMVDtgPktxUY1b0xd2QdAHxUNYzun0Ql9
8j394Qt1sCwfuEJ2oU/Fad4xMLv5FxrTMfJ6FjBhoxgT56SEJ0ljMP5snMRwx3M1iu0vSGF62fyP
WyQwWVBGbL/6CHcqA1q5YP2c+y8nv2MPWPTPgxu0YXsYYdgDm21asERNHKH+kF0sqDUkooWLRSbS
S1zca46tMcJIjNhhpwpxWr7MV0xTOVMgHeTau4ulgPtdwpw+13oTQ27wJHtzKYsdY2j2jual6xDA
mU0b1hsBbpSPmVP4qVdiWvH7nyf84Y7RC6tIFrEwKwP1F9DRCGQYQW/dmrtu7KUwYtD4Qp6FSh59
WDBsJjAWniQCcChyJ4CQcnxObPlv4SucytXKgKeN9au71y4x16RNPl+26EmHxUKGqiJSC/eF9/Tb
FGM6gGxRU7DjHwiaP64400dF6snfBCnKF/ASj/CzxJopVzI2/nDENuISylKg6qeNmxaateIcrqZX
F9fpmVm0OyJAp4uwb4NfUPV448evKRkrqyy+QH+Y3K7mML39Uro9ehrePZldHo8pJwBs3gUFEYVD
J42b9OODguLYlE5EXJKk88kj/PhV25CtczBxgEVOP+pEXoN9JqoO6FNuGD/zbGFcAR63AFJdniVf
CGhQ+aFeIbPE7oTxteUr+AXykdCpAGpIL43cpEo36meehYHazaPgv6ud3Jry2RbNwWpssImPpvnW
Y8F9+IRSDWl7o0mfZfEYg392FynFy8XG7g+2seo6g7LQou7NidmYWJQVukdf5WU065A0eqaoya1k
uLAwusL5ySPb41Os/PF20+E0xuFD+JrIlt130iu0wC2e0aTDj374T8YzQKZhY3byVMTIcAjzNjWP
A0GfnFLcK+W5/xwCJG9ZYAdOqjk0GOwsQgUC+fZ77541Vfvgt52Dzc3iVid3ufXQe504BzVwAh3z
n8BEWpZV9spFhW8VDe0WJ8nW4rTmsg69ft4azFeegK/0F8jxsccFoIAMi6UbpM3FEGFUlPMbqCIn
4uSQAB7+o/BplkIQcfdr+4HIznfQhILoIflZG3jaATNgNO8ZSXa2QLpeaOeZb66VLjE5sriy34Gx
ON4Z5Jbj4m+xwTpuam4HUAsdTeahDy2iz4ekbYMnv3yNnRfiHhtRLdQevyfmfYlR8e2RnbxpnOV3
+i+yOEIpMrRww1y8ywNmyf++y8XLhaDGKftHEkJr4EO0SW+V6TJ9Z0SirwRmI2d1T6WhrZ8GXRGQ
P2tranY3VsewGgmbs54SkoN6Hm5PSYMY+l6llf9lSKaZagXHnNGdMuLQgtLGA/dhyymCpnoEn6nI
nalQk+LJC66RSzR27bwKAMF3RX1ALleV4BHwK0k2icWvldPfE3W+huJ42vL03Ot/oMX/GiX315G0
qzcYCIBowaLr9wrf3PFnEaECgZxdPizL3f2jjwK2YviOrQ2EL6IA5aowYvNCGoGMEXEp+3RO4/xY
1odScukJ+uS/u3SdfEZLVW6DE57dpe+ZsGxUM+9sHGFDy3D68cQoxUd4p7hlIw7+kwBaPJ/NQtpP
HzKSgHpgG3gkSPDTzTeVOBBMM1g5FZGmOIOld6pKYLYXRb4jRzU5+XPMU1C/DJ8xn5yQBiJKUJs2
rFk5aIJwCS23i1vVxlUVbQXdqG9kOxvBe5OptMW8Cq6jvl9q5foHxPE946/4JCfNqtbuerYfos1T
g0bmn51X0OElW/r8kfFfYLomNVLqbdbU6pIBtkZ6lWxDY+cBlhGJa9zccMFfOITiLHU8aQ7409/m
Q0BgVXw7slzpNXyRb+QJtpUANHxtCVrhfNB3JOGYjkxfiGgKte3JvqARYnnUd6gIggw5BWgvu0AK
mI1SPYIhgTiyHVJHfD9k2TGSHa9ktmczVLg8PGJshA30jW0mWn6Bz1GPX001OS2wXrbVbxTWuvd+
p4g+ul7y0hOGJtFbb9tt6IEkdHpeUCKmBtMMTrLyAFjNiXGYI8fn23RI8dKVVXZjyfaOfTuPYFBY
kGUKrGXTz0Xrws+1nI3pdKTZfMuKFjzdgXRt/GCkVjKatNe6Uso04tf/sKnZg+HlLq86urSWSwjZ
tOhwvTDEsvktZHbkIqJ88KyiKWHCyfXa8RHCsHHjienNh25/099AxXJxH/SsswhgCt8P7BrV0LBO
4eBoml+2MgAZklspztaOLl3whRru0RnJAf25p0RPMtMhrOi1HprKXPs+jheGaraeDBlPj5GJozpf
eHK7KmMyr3ghgF4O0a9F+ZWSDt8pF+d+O54fYSlHHpPr+TpE6wnkxeqBains/gEVyKgee8Jm0ZWX
PCo8I5UFST/Tv2IG3evQROWk+u5WFzm3HNjawP1fvM67DU4PKAGS5diPgpZDaNpt0P+ANIPw9y50
mJeX661iVvy4TyhgqgHoZLu82yG6ZA9Dno5a1XQOSEeOG39KAdIkQS7xizOQzPiGPCBf6wVgvgMz
FgVJlykv9KIaKauf1HLXXfBGcaPbRoZJL1woz1iOfZyWKrsTk8zXuamivPvfRgjmSUIQfcJ0P6jl
5GJn7USNQB148rxFZILR+hCJJjOHssBFI6aLZLiEAvmsB8tBsk6iX3bWjnJgbasaQvo3Sx7z9mRs
whAWhG6O+yA+P4isDy8B1sgpD1WU4fZBQkUpPOCnl+86r8WP00AOBflPN709SUHEyF54VnxYKfTU
Bw+++8iZWxeB72pl07to3edhAkSQ3mrD7JKpFNqe39J+1/nHB7+qojPQsQPsEChEKKV/jxz1YZLM
JsldD6CBSxphQGzKwZMSMpEo+HRAOZ1+kYBU613w8YfWB1p5CLmLTt7LMyLwhPn+ORJaah6HWZSi
hDn2p7w5v0XdniLw2sIaz+TmZ84o3xhIBR1iLhqM73EtXPiNMT239zToUWRlX2/L/IG2iPyjzSOt
erXNYHRk+x5lbbDYr36tGWHXhO+3rr4mVU8v8n8zeKI5/TSj6iIK+XenJR6Uu5daH28c92id++63
zB804VG3WssclJeYEDjDsESqytFo+8HLwPNpOPTvVbKW3eCHH+qLyKch5u8h3/9tlVgI97M+4EKp
l7nOb1wSc5iaKdfucaubsT9didYhw228stNQVmud+5MJsH12I5+HslcP/uWAk+ULGD0qPMtjMrha
yObBxXQUcP04H/gXCff3tixfCabKgRoKk3Rc2UKlTUtdftYJau8ylNTM+BOUCIxHKskb8jDRVh+Q
gducyn53rHaojSFP+8+XKy3MS0u/v84N4mrZVuPmf18AYFNiXVKi29xnEx5hLPJKn9NM+BqTkjh6
TmiQ2dBWq4WWTy4AJLi5SVm9xaQej3FfIWneiIwL5ttad6Q9mDtL4ASL6vQlgYgWd1oTsdO3x03O
4paqzpZHWBFef0/ca/J6vLi7ra6cqQ6qCaZenCUaP4gmKJDaGCmRKd4cv/OA52dqzjlvqfUDEgJZ
h6/LHAs35ns8qk4cDPhlfhAmiGuHAaiAqTSZ4pbACLq4L4oIbHBZym5XBDuEJLArLLJOjPws+l3z
dvKaRAEk4c+kbEk6ICQGtaP/yZc0yZsLPSPN45trUdLPBzANcqudfe53u21qSXRTTO+SBKopkDa0
a9yHhIqent/bNw7lM0IrtK+cVgJImUIpFHMHTQdhVM3gMaZY52TrxFHWKdOjbDNIVexA6OA3hSs3
GfkrLA9okRZTO8xtpTL1Ria7ubQg2/o/GgbP5GmNFvwYbIUdd8U1WOZ0krLgBnTtxwAbhCWzlBHA
D54jBBVomsf5bjpVkhHNK2xVnK/1ocoIn7sOrzuKtyxmg9bqrLw8TgqucMeZ6zJevlTHwi9sVojO
JBH0m+sh1a0CdBlsC/gtPKI91bmoymX/cp2mC0fA901Pah4FzxzlXsl2Ymkdr19WsuzNkhrih6zy
goqys3BnDpOheg5P8DuuuBTSGouWxfVs4lPvtpKNYmsYOjj+5u+VAT91Yt5oXL7Ozq3S8KCChnvk
Nnt8hUYrTo01OJx0YikjMbNfP7x+wveXLs4LFLLy4UeUdhNiCthBZ0bsxtbYfQzYPJvmQKwydJcS
/RU3JEbB7ujVrzydixSOSYnX6CKJxMw3gtTOYVYvRoZX4GOiANGXC71oP0KcK6Y3vYveV3fl/FH9
2LNFJUfu4FGViEXALt1CAoeuXJ5WyL4wmlqCjjlh8Zmn8WbmXOUb4P0qujTa3KWr69tlGueJlKxq
dCAn2m5NYeaUKv1XqzcRWkjW0gO/DU4K1XNX6V05gQ60m49C+KpUWkmteWYj1w7vZgAaO9Rk8lqp
tF8Q6Y7klLkltYuY7yzPqm4md4IPx8M3T2RG9rMmEIqFNwv2jS5jfOOYRF7xCkP0w4neVZeueEqX
iNMEwdt1aK2U0GY9XfQBkK2YnAKxfQ21p85OB6sUuz9BufqsLIV0avY/WJpxypt79/cQkbnFuPPB
FEs3jcm6dixFcbDk6jxEO09G6Oxbzd3Ned8c2F3zIHKNd4PaWWIG5a/FoKSXraY8JWYyaI2Feknj
5MwihZirVCSkRfHo21cwX2+rEawko1FeBcl/LTPFvesoBE6LYQnrGhcjZxPQOsgfZ8/g8GtKUfDM
Mnyw7RJ+fotdMxylI+E1X8lDELUiOkroOVnNutTAdafMywMvoxRO774uwIkGM59ShcwvFR566OMe
QaoqCpqQhh2JIJiN+hsNID682KJjaDEmCMm5FuS46adURqVuGp35re+kbVJfCXrnyQx9t3zLckRx
xtcYiG+sDpzuikHQc/MjcSafcONUzgrS8f3Ffq4fvY87UIYhROie1Jiu0qY2rhzf7t/PU55+kWA0
6gJxVMBr/EwKoefGCEPdgdbAvXE/lh+y5jZcUWKYCiacxaUyymOMc8Wqv58SSblqROx0GZ/P3r/7
mYlg2xnrTwAtSkQE5BBpBPmQwQWMZU9/Cah+O1MsslQ+9N+MuSrc+kWYQwQqXjpsJLftodGRnYjQ
MFCOANBw05iA76JuYYnUlApC8032/43SlDDC1u4mtYbX0It3Bw693tQBY7f+0TJuNnEiyxTAedcE
2DPCx/wSfQS18M2xkItGOk/iWEg/8MpWMY1if9XuMgH78YeIUMlL0Fo0bzczFMgpsB4MoWg5qMV0
FCbgsLOgBenLLTcMxHaBbVP1NXftLc9gpLdlkrzUXv8k0o2yOIAzZVlNr+4JuWMy4Y5zZ9628BMo
wgrvhGWPBnGPAyhWODwWfXD8PG+K/UX+bPxRwPXv5rnTW17sf2uvdm/PJDOX13QVnshTIEvUDHTv
CRQmxyXWBGBI8WpHOJ8HZ2C0MGoYByXhITsfgd2rPnuryZisn6z+w664Lt3tLUBDeZmQtzXySdCN
u+dsQXi4ZNhatufYDXkP7E+PEkoxRUKoNcacHcND0Sk/5F12BoxZFaABk6FOHVAhn2AIWFem8taN
JrbCFPEdH8w7+5WUj6MQRa6f4KhaM41pR28JXQo4c0ZYemyI6OD2GJ2xNhBHMYhf578ZDR7QWHqb
h97Mir7qsJfPIVzTr+qBk3vRjM1tHme9/DUqwDsc9Bkv8hPliIYJNddzHlBLWXoL2J2MNChrI+f2
aWh83AAFjBYNCDQ1mhWl0L0bVeAztky9rl6tD4tqCTO7iLYSbP8ECbUo2zGMkFhY55ZxU0Hu1nkH
jU+8LnpT0m/rkzea+jyiWnT2AYcI6GFYs5D+5g4iZTy+L3YILfk30RE+k+zX5UMaQCu0+qeqyc8s
tVXWE8O8976KUssfBCwniCkKp79fKCMzrmp3Q6re9RThmBw3LtYudal5gSceykQ15YIQhpBbSysp
giEdGpNvwWKlJhCEdWt+C5vY+ud6IaCNv4GFQSiBFVr8AOmmoibixS2I3nYvIKY0+mxprV4Q9QSt
9rY/RLKQspTZFHMKNTEHYQewWYOgTeMoILHnBQi1SIm2csYiJo13grCuzM/whnC+I0JCqhsv1BZ6
TAnBAwCtMhp0E0GTJePQ4CNNhQE4dHe2ZEaB3pKP2EARfuqqSy9hECQZEiOswWv4jkrEfsuyhUQR
0lzpRJ75GLBMLDwL5DRKdHLwBtXR1vLnkNgePRgnR3jiy32Uck2FezqO+UvDhcWq9lhyh7RKN8Q0
mQP+08J1gNdL8g2weFIHetcHXxBa7cTw0PIkjOBwcNMuceKKkXI+EpainBoxPAOsgAT97voZFJ9U
X8HHUYM6E4GoK3W6N1f87u1i2LP6Ol89oUQOvub4bcNoYTrNWYzhNJwTNEjvmrNDFgZe7/TknptO
QWER45sal8CvcwfpRiPvGQWdfcnj9IGBTCijWzM+XNBlOc2Cx7nB3SIyv1No1EeLS674jebMzbYv
6ML3DyKxm30hSMM1smuZw5Fs4dSKNS2Er72NptW1mYa+x70NRXc3IWok+PPaQ12USz236D7nRRJp
es/V7SoyAP9lFHlzUfMxUPNzEf49nPO+HqiKea88uF9+YZI8yrGJvd6RrsvxR7c5sMZDAk+f3SWX
AWSiJ7QEYpEDYGCSAazgQQmbj3Q0BlG6h6SbIf0DcpBCPm+HUvrwjFsoJQCU3XQ1oBJduU9hWKRv
HuJ3BG3p5qrVUqejnrxVKGtbxT+Atqwz7LgRyjbKQgpZ2+4tpKPL2ccDpOx1J3UkdFjxYAa0YVnV
Eg5kqUx0fb2oqDnOgXadvupw+yoEgoThLiKxVpCTM+2DN6Bre5jVkMzaQcIjv0ReYIq0XiCXuCXa
8nsB0YhiUeyQKUQ9q39fTE0IgwS9I58heiMknze/WgAlyo6OdY9QXbhtXpuji7kCmLWdsUDqf8Hg
pt4kDLoSzdJsuqTHzBqF2XzliZ5MBFeRhNkrTJljQJ+BbCrVWWzb81wtYnxLg+ug3wSqRur+PhPK
clNxBePx+Y3C3dsbNWZpe6Z/QrLOjp9VYBCQBhqv1z4vhB6YQW7a2ZzAI8AdoaMH43EDAKDsANWq
CJHgwO0Tjr5YMCyoj+z/Enjuky4Yexon2rJVk4AJ5VRpCnqZrAu8CGA5RKDg/aiCfFuFnCIfS3p+
+1CWsfJAi7RiqU0hXFg0jQr9NqLuRKIzZjIBNdFrTPp1/Oid18gO5TNb6CfPKeyNzSy9PA45IH7F
aDE4+AchTFcNzuEPetz6oghyQGi6fGGG4tmuRwRG4Uhcb3FKke1lYt8Beb0uxI5+2cd8zJogmv3G
/icmid4g90bdouZJFjat82Qek8AGAbrkDz0h/q+LS50Z0NFgJk0ZNHF1qfqfq36TDBsxwK695wy9
pkmqE8ZQBGfc1Acjdma2m2Ple1jqvp0NSfTGoUrhAXr5qL6NemiF8oBmhb83rVO5s+9xSlmWzK0o
jGpBeO+4OO8JMownMrCBxkL8gsL4zQ2as7Wc1POdVv6T3Z5YuvQAN++ZcZ6qtpKPLKcSFUfAP6Ng
8dsbkkuukIi3iht1EYZmjvhkrqJVa2L6nkvCLahCjlio9ntABicXaZOraUKeDYDfUYYbYgdKx3cj
gijlr1A2hMrK0uZpKB3HHm8Pv8ZEfyfPqfDODMEh6GkUm2FeJSAy35Y0cAeM1KVWwHb4wA0MCgid
1i7YQFNhNIInIVdhBchLhe/jVDrRnCQADrCi+y9fkMctHt97zZ4s7V9WIi2wKBmljN2HCnBLi249
vqC1AkgpTcWowp/45R0NuOHLrLrtotLOeDIWSo0YuWydryK2aI3ETxCWyj+L891MVPMp0Fu/VnCQ
8ZlNHvSsy5Fm+fQtvBtABRW5X6vNB+iWyHnHumLjzYcqsi9iXDsYapq+6limpY6iWzvHMSer15Aj
OYk5flRqmODKJP1v/vlPewLm16Znkt46l4abkB73Gb8Tdd4sNuld2B/aKno7TwU3TUc8CLIfvnXj
DNNGgKG8HIxFEeeDE7mfLX3OiTT12wvDwilfRt3f34poIxxdoc9Q4REeTUFqQiePKMr1SXnv1KGF
yX5toqtEtYb1fFPyyf+rBIO22Gq8MjXq9J1aIewSK28u5vbgDw/QI0dBzUka8lVp0DYPkBaVgShG
NLx5QkNy/CM07iYu1GoFG3nTYZD6rmVXze+W/VfooDrX/szpuaUqKYfcqmPifanhf5NRrHDn6NGE
XWa5V/El8mF1wcMSo4auYr/RmN/CwlLe2djjQ+TQbH/gzn0uKSGi6AvAHCCsiLVdDBnMiaS/0UqZ
OaRiZtKSXZAkyiNtzp/0+wpToQiCaJiR4CDLjFmqnsKkDfcbchIO55wDYvoEEXOXg1zb0a7TDayD
WVmlL7cC58XEyYi2tm26SoBmJhYPWzZrEg41aExxFnH2C5mVhiPuUw2TsQW6OGpvshkAAdLp2fC1
sMT90zaCIDJsXbJ5MrVaOG2kl3sPgWM1gTtopSlOkLi5EXmNE6yvIeWuhiIUfS0HtmZAC+LqTz1M
1KdlBczrdwopy2lV9Q1JBs5munGDaGIfbpHCUU9PJk1FrwIjQ6RqenYw90SqB5xNrr6js2ImQ5rr
Pd2p8HEVwkezheys35f3aLS4I5S2U1mpbus/zXcNFfdrKEpdOrEbTv7HOtQ1S7dIIjIqQTrTjuXy
TKtZnhVmgBFQ4ML21l8nB4dTabF5UfsvpLCNmlfMbeAy56EwZoETmIEcrXOt9aVp3Xqnb4bIl5qW
KA6sHrKYUVqcMs8eUcD/8JF4CWkdPu1YIxr4kn6a3mYEbD9FKzoaJrEkPf+HXv5NtvHBAvWamsGL
9D3aWwSDor9nopVgWfenDw+03mxU/PtbxqRgFn9jXSOnUzzOFjxGisvh3RDZMDJHBxTwPfEE1eRo
GaFk/4XiVkSyePs9LrePu7GvJFdw4/GUfdFmS/gaSaR56lWV/JQIwt03uAC76a4bfcpADyKbckCX
iRfmBFyVjsCbS3mZDFwR3PeNd8VayRM+T1O9gyKzxcaq77OduR22j5m31c0JHey1AaI6Eli09jBF
J4gNapr1zhUpQ825u6kx710ha/PXysnDraYhVYvZFiexltMLjkSBp2f9pVjjgslzZa/4Z5AyL1lX
8xVlY6CHEffrHS/KLnX2b+EM5i4xRzC7cQt8Wi2hMc+cOdqCDGINmMr0HK6ooqac6b/LMRVJ0Ume
SLeEBCsXlpk9o9DEAhFqVHZNsPYh1Gz3hhSyz0QhWHbl4GB59IjvUnqh+8rjeMr97p8Ks2Cx/60o
vIxecnIDV8RZlQKognp1YnTJEoKxEG6mcIpMwrfebuFLhS3xC2tZN8JDoMzrhCWv+Qj/GjYId5vV
fIhPy+qT58MZfcTT2T9DezX1W5I5NPrrlWQq+uHTNCmhA0BrCVvotulbxQhj1vSKdwYVxznV2kt9
biOiJDwMDCqm1uYtvvPWw9lNvpOZna4BYLxQnCu6kWHdh0f8KP0J5BILR/495FCucInmtuaiNPHb
aAh/0Ztqjr4j+JQlmOCG8DDRZVmfCWLnsw09XRQE9kPgTpg/9SclCCtLENt08v+yjBY+1aJDotJC
Lu54MtAvBh/GiUSMClqvJolyX1iktIMB2Lu7MCGzGgEipI5HaSG9AsDFnAhwwY081vIDt9jJ6joP
neeERlVfn5xHoTOydYrzzY9Gw0QEwv/30A/JAWBdx/IY9GP9ziAXuJxjP1JlFmvN5A/7nUHSbS9S
L/pUpkzWl3/w8GW7zRAdweZL+9qPaB4/wvdA/u2FMpLc982l+z7mJ98C+xv/0pHSIfoLiiO7kWmE
5n5CsOjfx4Tl+CRnHE99MQamS8BNjNg4fGCLWUfuADihKyf2ZHo9WBmmxqYP0P1pKVFcF9gZ7YoC
OypZXaIyZZZmotOKZPcftS7Xm09ROVCSijhBHzxPGML6ltqcTLkzANBe2F9r0HtyERYGmdUoSRGZ
d6arsIi4nvMreYLbLtsTebyz1+zWjqemKIumerFLLYS8DuAEgNfsUgqtrQEPuhV2Sa5L5/6ZkE/l
byofGe3y5dr0NOFMe7HKQm5Lkqj/aM5dLFFI3Va1jPp98DnUPFX67al00P3w2Cfgz3EZs7H00dOz
qBVRiyVa8DezasQCNSiJS7f3GwgiXxBxBLJ+R6oVA9UAm99kdPYFIc9i/0PXGbPCncuVxHO5fiu5
bVcGAOTGMx5nG3B43DrZ2Dus5DDSNn0y7vkIurzv0hYEhkzv7rRcXxZ/DA2PQ3nXuJnycHvK9v5J
g0Dqz995aXnfc4JyUdQVsDq+Lfs33cOIFnNZKNgiC91uP366yQ2EyYNtuD97PKAVAqQuuSCGmiN+
g/HM+3bAiD5sFzqOWixTIU6yobUgLwywbrKXaxA7q1RcjnLeNvQOhmsRk6AIeE8dRmIbDpWdcmaQ
8fIZic0fEYv2PxHDRLYydVE/lGIp8ibCgldSo/+ib3eQXH8ED3FelkdU5sLLpOElkDH9ycKDggox
jH71GuVm+N0kBGuv3KCrS5D5FWnW138407vkSMT/tVZdANEMVs0idc41UeNkGkHs6QXqW0OdFG3C
9zcXg0/VMmQfSg+lwGkzgXWG+UNobaKgSCb6PqxPMEXRLNAHIyS9jCSOhVbduRfk1kEC6GiMS7WR
1wBq0Dhz/uGMF9lGuKVrYZIsu/zhsYRHrwQbtrmTDRx7JWOYJNY1L1ghulncAK9TTBeMbwaZ5j26
K1C5muIrjz0sFZohLI/ZetaTiNMw4f2uRQD1N9k7ks9+qBuGJRmvbPf51uFiEK/QFEuBIPy0E4+j
ICL24qWfFWS94SE+Kf1E9FCQk0KhiCbeZg1CUGQs88egVnz8amkNhYzvJ5WvjkgTw2OwjqqA0A0Y
FX5khkUkumfiyNbrbrDvMfGIjDMVbiD0la3bVZGF8TvTiFHhiqTJ6899kr9Wp+ZOEqxHtMacZg17
d9OB+axgyZFtf0bnCmfO1Z6sx27w4ei884PfwrmAzf8gLamP7i5JG3AsoWJlCAcqSo9YEuq+mCEQ
OBqI3Fd86YRO/RoPJBlukVP85YuE+8Rw5jD/cJQ9zIljkiEOLkBK29K7VlL9K68MKDstk3czOQ6z
JXpYNb2zQjJ380zE9oolxBWH1xM4PuwQ4W1QM6MuK9MPh/5sTpWwpxaAXlQc9P4+1bGZ5K61Jutw
qhHvLHddF1/o3ZOZbz2O4k+GM1XiU0fkk/umUBxji35CGpg1Gfp0gD4V9sS7IwRZmEddtM9H0TFq
0aWqKuCe4dYfegZweK6Igmpmdo42LRvN9CTsF9mE425Y5S6OGiOwsCAcm4wDCEOxv7I2QDLNtBWj
OeQ47sRF1jBUxnBbOiYR+Tu686lQHgfYLAAdOF66YIB4kSDHLY1N3Qc4JVfQ0nDyMFA9P7Tm7PcJ
lop4qDrO8ZaaZJK57YXl/3bmHynCbU3VImcpF0SJGLVQngRq2482MKY3DMssZlv0k5If8Tqp0K9U
N5vXFe593saaBqEzlq9VnwEq5cT1Ez3HnKDUAg3RWFX7qWD+O03SY7phSqrWQzRiuGVKkbEWYjhj
8IMKfvBcHMeeDUNr5Ms+lFNbr7e/6EOFdL7rYaJfbjxyn9nLCGdYTjm4V5YbtwOrP/vdEC27eoQV
mLBnmZvXGBDUHbwMawtbP82pb7Nl8YLR6kfTuwlxKwyXB29Cht6itF19/vYd2qcqn1V6TTgKqDUQ
4MmhmDIXg8CJ7Sjod33pogpy9f7x1OjwddoyZd5s2waf6y7o0OmM4uW4XWYgzdfA5uyVLs6fGZC+
9zZHcWLqtfAidED3jJS6MbWUI4Q99I8C9zYRKo/yUuxseJtmpXkG1WSfcgNSO4NGWsjYvF7jEnFw
kxz8AtPTb2QH+AuebiX3bAzNuqdF99jiySm+aOsu2hGqOLOHSlYTeGcv4KAJ8MiACwtfv1IIJDcA
5niwxyumRHxjjJEIKRSFo2L+geCjX/q3ChESZroD6BlBXpkhcbK5b2HPpqiCPVTv9mRk+Er9OrHv
oHFjVY5RtQAG8Ixiln0iaR6wg5wVyxnzsAeadoAHf6ME1klU2Qk1RJxVJnlVzhH7rtYnx9LyK/wx
HqQBICed4ZmCZT4d5le//8StQpnehPiaoLuIne25ifAp03x6qzVWf05AF5YwmBtJdf0xUshDeRrM
XVBHiOYgq+EPx+FBWEXFh845FLaf6YslTuOeaNs5lzb9JL2qHDHDI6sq7KZsrZ5RPlW6u+rSp6c6
R0qzyaSHUiqL4G4sHdcYEBC0byOU54TOmt4oXxjr4ugVUd8vy5dYo+YOD3f6qc4z1a1meR5tzkpn
i8GspN5c0y6SgweJGkJ1ZUWIhABAekIwRqGSjYNCibc+vhLsr8OEVUUbABi1vjDQv7T0Jank9UOA
e53ZtpDfSX8oWKd31l2gEVFVHYFL8os3A6wL5uT8KtT/xIUIyCp5BoopADXSaqklJRh0cuDMJPv8
BMRNWKnByeQdAM+XKJLeX2ZIhSqbmWzMreVe7a6STFbo3LHEdbecAT7dS9aUwa1Tg9gEC6UATCJI
XuXSbr59mlckunPJNaljdIBj7afoWa7J0rpH/4Skbo+zkX5/S3O5YJNLZLBfKqoehejJl7m/EfL7
AyDuAbHv4QjkZ7RJdD2mJtnkrLXr5MuhmoZnYdT4wBeLUI/D3/ZBcw+jsXYKbc3PCba7tbPx1nrH
Cxq94dr0nOfLIIChDwOMiZ7guuhoifSxMyzxZwTyhsokIs+StcIW/2x13Rx4RA5dMiHI71aHgFDp
mfB+M/w6wi7+rIu712ONf4tbmIwbiuJ/VAnr05bYRPBHUA5WSt6Kofss3F0uDcBkfeLSl51++v/4
vT6eCRkCvMbPfxRCK6QLHOLjX/aVdiiq+JVRCKfyWHkV/zN024pPppYtFGdrcew2Uwrhe0kQPzxL
a/whmmfwtlOJ6IremnPYE9hR9fVemd/bWKGz1gFeYsT40c0nWjQZJMi5G0vU4/SHKJ/N0gWQu1sy
e7EYwzH7Y1zAPCJ4k3FiFX2X8BKV4bv77klNCMD/HdAHAEEMfM9virxcT/Br3rfzywb+249PYeBn
L/0spgt/Zfw0qRzOOP9IdLuht41n9opkNGlpQNXnWXp55lBF3xULpUYmH2Pv4HoizgbjtIxoQt9X
u/iiu7LX8xq4JBdmWGOKxLtY3z1YXrBwpKTbFLMWY30YrMsPnIRgenXXXiPm8cZ9IYfCNmZA//7f
uSxG6atEbbptf9/uXL8XFZ9VMKlsDViiDct+b5rNNuKKssapZdISmPt/SaDdJA6hNU/dMtjWvdFk
uRnPnTLkgDx9MEnk5e8erFQDth1l71DXKIRkemb49Bdo4o5PaGDUKgRSpZ8IlMkD6snoTgfmZ2w5
KesT/XnjioGBr+421xWHCwOqD4Cl+mgJQpHpWM3qAa55kCEPn+2hjCDLKwoW1cWxSGc0ghiKQ1DU
kXUlpBGFw9cgfV/Utw2b6+fr09ADlfzK9bXQeHwQ2g7y8tLJU7IzaK1tuHxRf68u6vQPC453Ke3d
IeNglz/T8mnFU6uoJIshJxtDO3kTytGFiot6giscLGll9nirOCrKD7T5rdqv1jVv8ArWGhL6Ithu
7Po/YMrx19g4P7B6lIgE8FuljuRX5FkZM37+13fMYLTl6cYX3n2TMQR7vbxsQMrVw+npEZZuaCjL
Eq8e1PpyVHjQ6D3ThaQy/81jL5HFdr55c1sRlmVkjO2tcXIkzbkdZEn+vElUlhohXhnkTja64fn1
/h3y452ah5HlM2oAdMG9vnhV99m2ZciQqwf8RtKxCU3wUWajp+MpDohj99G91z3o9NejsHOJ75qF
ySmshsZztK+Go5ZWpOiwWpELnfkdN0Wgx3OLfnUqm4BIpdIgUuOuVK8MpuG5e4SDYK5fe9JBE/8C
fsF2yzwG5YjuwCUkAWgCWcnGUXD5vQnwan5loR54okhiBR1LBWcQpwQuUpuZEdB1H282A/acZwXf
6eLIIPLY7RZlgxWWD6MaESbtCgXhKXR0bndOyoIe0wraybUupoCfJq+6ZRW5/+kbq9Jc/j0zcK0+
mRVhEOEljasA5YW5KTA8TZgH66Alx7+UwP6zqeiYs8lbY3lTLuc9SV+VWqHqwFxEBna0vM0/gLkW
Vq4rcEYFrXvkDuZwOw4OpJamonkT7R79Z+eC1wqyzE1DFmwl0RC5R+obXWdIxILBw2sgNGX6x/6s
ZsydG3FhlSSi61SpWLM6cThRyKlF2TqansRqgiuQLkq3JwrQ+jl9XRfc+XiyJe77X1uohdux05eF
MmpN/APaVi9qg8DaWTF3zCDj1SnTMCsGMzhd9axd/YHKuE0l5SZzlCEI2aZsgOfgT0xpqclsGmuf
aptr8l9waFbIe33LmT7erCm6gFxLA2tZMMIuyNtYcSkNHGms+XMeBCE0dKFRJY7Y09U/FAMaY60q
bxnOQGyA2QQTZItXleplsr46aWSzKcA79HkhhsyuiNag/p7dT/3yYTApPqFk79maEAGSQjFH3QTr
mufmXmsgLjuvZE+9tIK7eTsJ/ML+e38h8BamwkN37wrvzEA6PnXZRdb3HhkxqtZN35CEWq2LsKrS
BgZq1Qyn/6ItrC4MQWI3bb35TLelkGjCS//GpGQQet1SIQDc8ocTpo9dta1xNIOT7Z/AWXahe6IQ
4DUb2YKqFjKEv+FyzBrf043H8PgNObfXKoMih050RvazV/7hRGS+g4ZaNYQlre8a3qd0nCs3JPtp
mhPYJCZ2qpzLltGFZ0/EJf7JdpqPFkKJzA6+oQLTeKRV3hp/VZ+LiscK7/l2nTlvmQg5MIx89YTR
OoouCeBmkxi5V3qlg91Br8nPuPJ6zOnX/kbeG8uuBDdsgiVTCGApfhxL5CI1IPJ8hDKGFdwIMJox
5JVlamq9RwLb+XYMOmrVNOJOjwbfD8PM+oqA4xmWFZOlFg3l+7HWmhExbMjdZoHZiLbbbTWegltD
WWoTranTd+oTz8vnP/XMP87Flojoxi0NdxOPgJb8yIFPnIa4Ecpwlys30Sd6mj4Ko4deeu71KxJR
79OH+XUfMw9rC8S5htnFK2yWTis0+0gBZCYBN6qjw81cbSij8VdpZ/2kBzrqvtM3NcLDPP/ypMv2
JFwI/JUZfjeA5Qw7yen7K1NfoZ5F9ANOXQ6tN1HRmCSIxtZ4W04XXzk5iAR10b0jUBO8jBzB6Qky
t6N9/kLhOTY3vdng4I9wRCZbP4TT2e8vzxh0FGAHg5umxxj7wvzVmTgjfzrxH3rc90FFFlCIajKl
Xt1NthurP9V/f81FdvSxo82PfQwMBzqM/Gb7yM3HPfvKfUikXWJxLs+STqYEDkFssqm1g1hk4hNs
jZecHM7+ju/VAexeHs4SySXCO3nxMULfgu4KAAyOcV2HEIpTwJuSUYvK/yjfi6RiRBb+mX1vEn75
9sBLS3cCiMS2t1AgG8mFRasD/SEojely0lL/ca8D+XrzlM2OtTpJrtHO8fAV2SvrRTwFARcEKaKg
ypSrgPa6Xc9AFxMd7eR49yx0SC+3pRBNQvmgQ9+Gr1yijKtx1P58BJ4CnC4kHS+iyztzpiFFjuhZ
CVnN7MD4OaBnG5FKM3hzP45GxkZiKHc+yT3GuNeMt8XORc9SxBWc42SD4bwSa8SO+nuSrhMf2iqJ
2L2aGuW3z6GXpEqnOspg2iehEGhHMtSsksT2RGjYFp3Sw7jOS2ZWTBjB4JdB4jDb4D09k2gZAGsF
nPWiLbyOyHq8v+NxqpG5hkJMPLGFjvIFG4NaSfqOiviEsDcjsq0UNJzQdeTJfJZvF8xWVVG3jUbY
IR9xEGQkUMsAci7y2fabUtprrObzUfFiRXw1KABVR6kJiPLGKgb5ThxZ4g3EK1PRp9QWwiOGA059
spfgr4B7K1hfr/uO4fIptQK4kyJ0t3p0f25Q9uL30CYdlPnPvWvlQ926/q6yOBeECHOaNNC87uFB
dVSyXADPFpCFH3UcW2docBOD84t3HopP+R9aM7brJw21h9X3+s6gkGseoMJh8+3+rWD0kzPBlE3l
9u1u4FLJ0FPwGCgDoEyydfn5lts3oHmZYlijl/Zq7krzGfqIZpwWLHz8rWx3oeuLdHVhnz9Obth4
KnDQT2PtkvdzIi36bot6iANgqXENv2sYzKJ/G6szHkSFGncXH3/ncqA+faVkKGipsPC9u6rzk4Id
NlVdoi3Aru2f/G7T5mKNSVNrnPAjBEvrAsviWuE4D7lxek0TiDZga5NXpqGA27m0n5+VATxv4fCk
+qw/Qz0vanmFgvT33SF3Nx7Ic3RKZoNVq3jgggtj6kYveip/hxFtWyQ7+jRY2XYdEfrGlJZ/gfKx
LIw2bp1u8pdZUZaBHPObf0jSTrcDXXMM9QO2p8R8nj93skh8rvNyHAdO/2uxh0HRDeZ9EGqHcbVl
ecYzozEvXi3VWwwom1JWenHkhEvGRiBMvDNnPn1w6tNulLOY90nmzt9qidUASmFqNyMeTfqnETCL
OxZ9AguQq9DtkC4RrssNoW0NHPS9nIJIoknEQf4cY9DSD0CTYvkRsXgv9RkXLJJBKpIoD08hUCjO
QlBOx6Dq0maY0a5Dm3yJtOfQeltsFpNMtxmEE4GZOkIfGk0xJ6zYtHEsQe5i96tKf+GvP1B+36pz
9LPELEiQtOeMDdwzmU3jxm6IYYjWhWK+Z1bbDZfny3cWbAeTgc8nBQGmnwXLNUtnGYF0HmgTuOvd
tKTDdY/jmRaOzxBNmoYHlgRvG3Pj5QSvP9kvFDJoRp0H3UkNLvZYGOppRAISe2sBzcXvI5VaNIgm
Xk5XptfeudfNe8JMT3+KH5GKWlAJDIw+k6iFGpP7YXWkDxRRrvIPqX3B6c/VG4n9AwM1cRxC1tYt
s/FNfTY/d8HdmMsw0Ixc+O4LUaAjkWvMAslEuMhonIhdnM+EyddQp0/vb0bFO7gk9jmc0ytjke8x
b6vrdiOFoapjUO8g+sGEkaWqIFm1BX0m6h1fKXaHKTrI1q7JDZYa2VKitbKgnUoow6qyXEWsmIBR
nSPy7mHd/eaAP0pBZFwdnoh6ydnHGGWI7Ud081orCZv1Ffm+9r7QcxfYzMmT6msys2CTcXoL0WIc
5xeWon6mleFRmmr5WGLTxHdgpGY3tpbECw+HRLYiwWbIxXiwJGhqri+rHKOyEaZxGYkd2NbQCsGX
UT+a6vF5tga1oWUHzKXpsWWAH00vROpybacw3WTHAJzg/zj/Q4zF2JRvvav8dVDqsAfcSiDLRJ1F
WAkI34D5WLhQFY34GSmY4BBhpGJDZcLjeQOGL0QCzE/pLHWZKL3cKeO7rQCUB08rCJSlUW6/pcwa
bQDR6bb84rWsylFyzHu/odjyGdk7D+zm71GZUaH5KQkFNYnaSEv4bzMKtDpE8a4ldze65A7T3YO7
GL5Jk2MTToDDrtzllJnJlTbcBKZACxgUoSoia0IBY4X2VE/yBkWnSw/2XGKxi3Y2Wlinlu49ovT4
pU34IKNVpgaENhYG0Qq7NHkWBI+Qb1lQhKHautDmuKgFPzonaWEb3CHYSEjLWeyqR3BVoMDnInhr
x/acFHD5Vw4zCf5cxTGItcrej6L836oXhLdBPB3MJtYkXzQkroWqGSEL5oD0kY6YqT/FDSN6eIQ2
JmxsYst3NJMJ/XxZGZubN9YbYMN/5kCvpDUfPJzsJGf02Ei6ZjUJPKsmYVyN6JRiVAYbJaB3YmWN
JNJ4PQHwXZI9ucc7UsfXTBNNSBZq+bDp3E5jXwFpSPosqBYpY3cYqbgvYBZHxYT4/iuaUZtGGdYK
GUX3QE3Sef4joeUGQUO9MhuiwCMO6/3FEx6roE79WxPgHUI3vb5jsusGV+XluujHoQT5Tn0h+2tj
I2L5OIcvyzy4S6GN5U+dz1tziB1K+tZt74qOwxj37K1xoQlZ2R3QPkHU6PQ1MKn6nL+7QMV6P5g6
zpFuTaZkLiGDgdy6Scjb1/jlP60bgmS4BRqG4tBLi9FZaGp/UDyOfbh07pglu0Rt8QpffN76cJP9
og1CztaWVKWG3NQv8ssTJu12YJATllNoOFju/zkCGX6JRvrSSj8EDnRFqvrLLx/6JydXobCw3pnw
Ez9KaG8oYSU24DMJa/9pC9WSwVNP29CrX25ZaWUwrGm4iEhAf+R2qRHNyCRsD6kQDq5TSU0n8tsV
XdNV5jCmIomKLqwj23yd4QG8TdEJPJeRN31th2qQ7avPlMmukWIWC0VM/TbVmlHiScWRw92sTGqB
l7haTh4Y5IOw7JXnouuj0YlQa6fz6mXyeovqDtYzNdY8FxEDuiWKscW0KvrgW+BTdkSRLs3MSF/g
nrYAg4b4tacJDL40d/zZUPPzMLAi2nW5aOlZ1Y9HUUPEnE3oUwzutuIo4STsXB6ubCsATEEhhYRA
NvWctTIMHWJSmF58e32rizxnQLRQEJNcM9wJ1vMDbAIj/I/bftLwz+rFuxFCkj3e0HI41JKXn1fq
rR/Wt4UHYH0wERANQlDM2/LTPAc46JowRtjPh48JsemLai8QAEaxn8OtE239akcJs2kVjDm1DreO
W88gqhBdUp+RPd8Xs2zvCLII/2FuIz1mV5kj8j1ZlLAsMlnPWfeKeZqACbSVKw6l+j6nwPJXRwJI
7TEZ5G5ae1LI4nbcc4hyugzhSOPYpV1KGkuT+kYXjj3PaY/0wKJO5RM+5e1iQkv/wPFPxNYDQaAe
bEBybDO6rUlaEav1YlV/Q1E4Lo/Zqai/1syv9LFl3TnTOBv73cBFS6Xlnr6h25VbLEDkcZnWxRDo
90NS4JPNXDwi+9uqcF13oxqKGBlbsKk1cjEU5p4CnW8GBHsKtnqOEorbPhBBly+Wh420gvA5BHSj
pg+OAfmcOGKSlQTImSS/aTFCpe70MnCWHIKHo1Heyo39nth/sbqAfmUVJsuWkLgqQrvFsUSQLRGI
eVvcooBUVg+5Xkcw9audUR7uYxohUBFBq3OOMZLMj+yZwWkBbN2HvOovqX4+UUT8JrXo5EyIqIJ0
hz5b4xUKp/UZPPAAbFqkPbBOxUforGhpZQmTgn9GPQRwUIDVTy+uyOxFx0kf8kSpaWcRP4/xVVrr
5d9KDnCkxqWC3c2jOPXyTgRH8+0oFa1LuymwzuKanGQRcmyEQuyaS58QHap0kxUraahPgQRh7lGt
ewvhdO9p77KJApy55V9lhB7Y0InWxDsbWulSXhtlL0GLMYX2CMA56vyOj5vFw6cGRvLlJ3/LRhOF
qus7l9xRf04BOVyPp/8lNbBmmb9a9vthM3w/VQUQrYRNoASuxJf/g7qE0v+cZfd11vBiQVKIszyS
g8QHuK6zT1gG0Kw6ZyzhGZTJxHayCJkR+ikNz8qlJ19szGHDOxE3hwIyvo2hBNpjxEUz7czA85ZZ
MrHjJofZA1mJE1BDetC2kfbWebuFXGE+p53RDsW1OPZLRy/nyJFuz/0kOGFuQMwL69omaCt0yK3e
t3zIFwnsHNhK6+h1+s/IdcjiiNuxrQ/lml+WAVktLUWSt/VI3uXJnZlEO0czJgw9ii5mRFHeY9qw
ZbX5x3XcOrWG5upOqDAlnB8ivYb0NmkOx9xe8IvXsr7EcMXdpTR30Fmqh0V3sfd9+1c1RHvjTxSG
lszq0ajFQpqBspkkRwI6hVHGMESzklr01TyGkupqkLwXhZd1Sq+eDwpUHyj80KdMqDX1L5kdNtW3
D+KVpYlp7dt/E5qH9WmOe3MWqBOzVo9fMR0jmjzvJpH9UCNABBvUszrkRO7zDfQVIa4ZvOOOxqgR
iD/RYAigWvrGH9Ev3U+roOYeEwvMCHZp6vGlzNeng4ZcAsTgpgl8A0WG6OkRb/s1LNGcR02shcM+
viH8mVYx/h1tQaZ6HD7GqX3y1zbjXiHiNQahbcf6TxQFukW3ppkktdbk3FxfHc2as4h5uKx2QqPm
QkbrjWLGSlUk3u9bgE3Zf8W8OWt9abMHKmQPTc8oN3LGkIj5s685/qyEl3k+sGx4BSOa8Gzn5ljB
q+9gmKcGZXYYare8/fmknGnHPSq0AzmRwM3e8GDKQZ9mRpydPhnzE2CL3XUwoPaYTi79oaM0g6Zc
BHquYZ8yyC+MZ0YQBWfPRkzx6VgTEZwKzrTD0t4b32SVCfTPukoMEUdviax8MHDkK2Hshm6j11cK
+dnmd8aHvMDlZeRCZG4h+7HuqoeREAyT+sK0//WQdcRrZ6aswHLASW0pIm+mtCMU/lawwMtXJPjJ
EViSptqoWebS2Z5pDRZeuT8k8CmRQF0HkAt9/Vz8i5ZNP4mpjPmOQihZu4PqFlJgy77pgb1jwyIZ
1jgXGPo2P7Dh5p6tVwl9I5RdjLaMp3mpuNhypm62M0V2gDhfsFI0RErT2wZLyzrKxa2/qtZ14BBw
EWSwqxF5cXw6FbcrwOlVkh1e5h9Zqevh3ktR/xLXajxFOPN1kcvzzORuF/xsaQ80M4N8W3CYY/VC
rwObjy/EaD2Og5evIivdj+wIg5ZNdxezp2ILx7LxssNdfCQi4CoDlUtzmcvPt9+YKSvSOywfcaRg
ZmOqX+m6ucn3Pnfmv7aUNl8FSwXf42XV9B38UkYCfZqb2hzmFUwOAMBge7fdDNi7P+3xE9W2yhIh
xrBgGeACpQEdj5os85vAyyI2A7dCVTSHSA2kIyFNPB6bPAGFDYc/xOfSf+DIFs9yxErVq/v4/xbZ
TbysI27RchNux7DNPF3fvYLZZHHepsSMJZnJMea920cJo/Obg5TcCtxVvVRL4MKmqfruXbItTMq1
9EIe/Yw0X7feZ8ueYTYs3PItQoc3Q21Y8CxOh9nbeovdK2a4Lcm5cSoD2j1Xls93qkNo2sTNGGAM
wZURmlgY/grXT8n9Lljk88OIpD/HGh1C4CaiiEcD7qQQ2XvRGGiV3KFdSK2zPUzTOlH8uzfqq5A8
ZUGsHe6UgxRbS3Hejxi+1XWzSTZwAChqUjuCu35LYds7oJ0GgEgr5nf5k1Au4+RggtaDE99p2Txc
j/qiHQEtMVkdRMT+z8VFeRKpQoDnIeC9G5gDzsLWBlt/Bbtx+kYhv4kFFVdLqmqVoZz1FT+ovWu+
nFyLt3+1OEHuEzHOsqXrcgDujrnzd/iSrsPr4f1dO3QwjIB3TsaS3sCP5xFjaAuaZc0FRWftHLB4
PA0Hlm/eUIUqUQFb16PRRO1w6sx9ajkm7xknUBb/kAYeN3kQKoKhnWMuynW90hZKdGeYq7Lrh1iw
F+3Yk75gKp3ymynQvUCpwd6kkC+O+47igeGNu6mMhh4Rj9gDXcJ3/Z/IG1jpHpH35C4enMu73+hA
SSHGfa170ykdHHq71mHMgs4SbC5C1HHPJ0jxxwdgWSzQ+4ww/RkFinNf07eTl+z0rDf2j6h0wSLa
ShQ2zm4QdDA1dfbAi5XuyikxYmmc5tI8A4Qawfb34zshPBcu1+KDw6JI1i7o7bAP6Ze6GFBQmjlw
jPUs8WgtkGbzDhHVrUt5oP+NuPUQXwAPxysNF1yN7ZEE8CN26apMGMnmD0z4F9MAW3h5GMkODclv
7Z5ihFLUiT4b0bTMUt1TIUxEhhu6tbdWPM3IbSAwNo5e4ulSU2f1/V8c7lMKM2XPQ3s4/0KDyIQ8
ZzIBdmrZdNGwR73zS8kRv47wx/jcCPSjQ8uhccfrGug0QYqPxDxOoWm8Zk6q+Ajh4Zn/1j1/0b6w
/YhpRLQ/Hm5cjWo+Tg1/3yl58iTyFayoyT2K8YdrXUcIjS9hNi/Q/Y7HiNxqWcrgrBsd2Le3yFhE
vVglMRduy71BSN8bO/0pa3bAcetzn8AjtgA4Vc3y5qHt5OdoJficJg/GroDqG+aQnLjtPEtk2PnX
yWRS6ZGuV2+yC3Tjak80YXeOEPSgyTwCKNM+jtpdyrHHkS2BlAWG9nRcmH10dAK/TosjVxV5+0SY
7sB0MlsoEFHL3eYESXrF/A79ElkGUuwxEgnGGuJclkIfVPgynXeEfomzMQaO3FLJv2abLHs8E3W3
W5HBBzYO8aa8EFdwEBMQcn6PLNViBee/nqUxhiR/sMOQoFqxULv5siJi+kQJB87Eiq9RSH1/7NqW
cVgBnPywUuUhn5lf9vWId+gm7dglQK8sSpXGjZLJPCdjnBeH9UhX1+AHGJ55AnPHD9TAwpvKdZlE
uTySbWATu+4JTcq4tjVQ6j6cohwZ4dTPOFBfn/6SzLks5eXhaLpi/i6lLBdBCPA33Vhb2reMFPkz
n99sDTe0kh8ZVR/9GtBaEeZxrliWbifYmm9DLOpHFD3imhnBJ2ikrasAbg/5zxNG8tqquIQOR9DU
feV4DOrbVGPM0XPepNx4PBiKyFWM4KSH2q8nOHSuwKVSy5yUNPRn7XodaqjothB51pdzryC9DeZQ
DTZiqF5IhyblQrEDQaJ8mMNl2v8UUETB/95J0UTYDc6ANf+AQmCC2JRv81l4G+iTn4baVnTeP25G
nsl/mAEhTiOm8pqTxCoF3NWp38Qq6TNG0lEh6S2eg5XcUn5ZkjDCK11Fk9Ioz9L9oR8JgGU06PLv
pz17A1SJZVLuEV+1L2VT4Mn/S4t271mdX/CUPO2HbI1DyZSNVSnxNm4GFJxB5qfOknyMYEQbZ6V1
37tZDdY9S6/MOJtmdi4V4d1owLr60GEBrNM9v0CTsDoWQKSaVKcTz/sd9kf2aWJhjjxuLQEVPZ3t
03WdEm0Nt6GCa2oogebZ/gZnLvb8WRKq0D37GuYlEnGOs7nFpDJlEQF8awWj878U+GkICwJ8nJEr
WdVOPT4EMH4PIg1ZvT6QMlfDM2jwDpTSrJVTs0zZF+1hgBIZceijfUL7ed5FL2Amsr3wdxnxArHw
HxzhHuPtB2L3K6cbFWorBzcrzjx1J/olxl18yxZKTSuYTzjTEO+lxf4oXPfsR7+fMxReR7/wBSOA
ndc6wrbt+iHsJ5YI40VCFhIbnAV94N8DgxRNJiFVLXGnlNFhvNp3fRsX29PD+ev8TxbbQgpVUpxk
FC8ZyI720KFJQ5HVLjh6cM+Kf2Hl8Ca0GixO4TtPbAi9Guatr1J8X4ujUAYCosbwdIXgbMIBq4TH
VE60qROlcO2anHvhZzWSBXmIuQbICjODyJra4hrjDksH/4W6adJEWUxn3JVVuDOA
`protect end_protected
